magic
tech sky130A
timestamp 1614098583
<< nwell >>
rect -85 385 200 1445
<< nmos >>
rect -15 1730 0 1830
rect 50 1730 65 1830
rect -15 1480 0 1580
rect 50 1480 65 1580
rect 50 250 65 350
rect 115 250 130 350
rect 50 5 65 105
rect 115 5 130 105
<< pmos >>
rect -15 1315 0 1415
rect 50 1315 65 1415
rect -15 1065 0 1165
rect 50 1065 65 1165
rect 50 655 65 755
rect 115 655 130 755
rect 50 405 65 505
rect 115 405 130 505
<< ndiff >>
rect -65 1815 -15 1830
rect -65 1745 -50 1815
rect -30 1745 -15 1815
rect -65 1730 -15 1745
rect 0 1815 50 1830
rect 0 1745 15 1815
rect 35 1745 50 1815
rect 0 1730 50 1745
rect 65 1815 115 1830
rect 65 1745 80 1815
rect 100 1745 115 1815
rect 65 1730 115 1745
rect -65 1565 -15 1580
rect -65 1495 -50 1565
rect -30 1495 -15 1565
rect -65 1480 -15 1495
rect 0 1565 50 1580
rect 0 1495 15 1565
rect 35 1495 50 1565
rect 0 1480 50 1495
rect 65 1565 115 1580
rect 65 1495 80 1565
rect 100 1495 115 1565
rect 65 1480 115 1495
rect 0 335 50 350
rect 0 265 15 335
rect 35 265 50 335
rect 0 250 50 265
rect 65 335 115 350
rect 65 265 80 335
rect 100 265 115 335
rect 65 250 115 265
rect 130 335 180 350
rect 130 265 145 335
rect 165 265 180 335
rect 130 250 180 265
rect 0 90 50 105
rect 0 20 15 90
rect 35 20 50 90
rect 0 5 50 20
rect 65 90 115 105
rect 65 20 80 90
rect 100 20 115 90
rect 65 5 115 20
rect 130 90 180 105
rect 130 20 145 90
rect 165 20 180 90
rect 130 5 180 20
<< pdiff >>
rect -65 1400 -15 1415
rect -65 1330 -50 1400
rect -30 1330 -15 1400
rect -65 1315 -15 1330
rect 0 1400 50 1415
rect 0 1330 15 1400
rect 35 1330 50 1400
rect 0 1315 50 1330
rect 65 1400 115 1415
rect 65 1330 80 1400
rect 100 1330 115 1400
rect 65 1315 115 1330
rect -65 1150 -15 1165
rect -65 1080 -50 1150
rect -30 1080 -15 1150
rect -65 1065 -15 1080
rect 0 1150 50 1165
rect 0 1080 15 1150
rect 35 1080 50 1150
rect 0 1065 50 1080
rect 65 1150 115 1165
rect 65 1080 80 1150
rect 100 1080 115 1150
rect 65 1065 115 1080
rect 0 740 50 755
rect 0 670 15 740
rect 35 670 50 740
rect 0 655 50 670
rect 65 740 115 755
rect 65 670 80 740
rect 100 670 115 740
rect 65 655 115 670
rect 130 740 180 755
rect 130 670 145 740
rect 165 670 180 740
rect 130 655 180 670
rect 0 490 50 505
rect 0 420 15 490
rect 35 420 50 490
rect 0 405 50 420
rect 65 490 115 505
rect 65 420 80 490
rect 100 420 115 490
rect 65 405 115 420
rect 130 490 180 505
rect 130 420 145 490
rect 165 420 180 490
rect 130 405 180 420
<< ndiffc >>
rect -50 1745 -30 1815
rect 15 1745 35 1815
rect 80 1745 100 1815
rect -50 1495 -30 1565
rect 15 1495 35 1565
rect 80 1495 100 1565
rect 15 265 35 335
rect 80 265 100 335
rect 145 265 165 335
rect 15 20 35 90
rect 80 20 100 90
rect 145 20 165 90
<< pdiffc >>
rect -50 1330 -30 1400
rect 15 1330 35 1400
rect 80 1330 100 1400
rect -50 1080 -30 1150
rect 15 1080 35 1150
rect 80 1080 100 1150
rect 15 670 35 740
rect 80 670 100 740
rect 145 670 165 740
rect 15 420 35 490
rect 80 420 100 490
rect 145 420 165 490
<< psubdiff >>
rect 145 1815 195 1830
rect 145 1745 160 1815
rect 180 1745 195 1815
rect 145 1730 195 1745
rect -80 85 -30 105
rect -80 25 -65 85
rect -45 25 -30 85
rect -80 5 -30 25
<< nsubdiff >>
rect 35 870 85 890
rect 35 810 50 870
rect 70 810 85 870
rect 35 790 85 810
<< psubdiffcont >>
rect 160 1745 180 1815
rect -65 25 -45 85
<< nsubdiffcont >>
rect 50 810 70 870
<< poly >>
rect -15 1830 0 1845
rect 50 1830 65 1845
rect -15 1715 0 1730
rect -20 1700 0 1715
rect 50 1720 65 1730
rect 50 1705 100 1720
rect -20 1610 -5 1700
rect 20 1670 60 1680
rect 20 1650 30 1670
rect 50 1650 60 1670
rect 20 1640 60 1650
rect 85 1665 100 1705
rect 85 1655 125 1665
rect -20 1595 0 1610
rect -15 1580 0 1595
rect 40 1605 55 1640
rect 85 1635 95 1655
rect 115 1635 125 1655
rect 85 1625 125 1635
rect 40 1590 65 1605
rect 50 1580 65 1590
rect -15 1415 0 1480
rect 50 1415 65 1480
rect -15 1305 0 1315
rect -50 1290 0 1305
rect -50 1190 -35 1290
rect 50 1275 65 1315
rect 15 1260 65 1275
rect 15 1255 30 1260
rect -10 1245 30 1255
rect -10 1225 0 1245
rect 20 1225 30 1245
rect -10 1215 30 1225
rect 55 1225 95 1235
rect 55 1205 65 1225
rect 85 1205 95 1225
rect 55 1195 95 1205
rect -50 1175 0 1190
rect -15 1165 0 1175
rect 50 1180 70 1195
rect 50 1165 65 1180
rect -15 1055 0 1065
rect -60 1040 0 1055
rect -60 780 -45 1040
rect 50 975 65 1065
rect 40 965 80 975
rect 40 945 50 965
rect 70 945 80 965
rect 40 935 80 945
rect 100 800 140 810
rect 100 780 110 800
rect 130 780 140 800
rect -60 765 65 780
rect 100 770 140 780
rect 50 755 65 765
rect 115 755 130 770
rect 50 640 65 655
rect 45 625 65 640
rect 115 645 130 655
rect 115 630 165 645
rect 45 535 60 625
rect 85 595 125 605
rect 85 575 95 595
rect 115 575 125 595
rect 85 565 125 575
rect 150 590 165 630
rect 150 580 190 590
rect 45 520 65 535
rect 50 505 65 520
rect 105 530 120 565
rect 150 560 160 580
rect 180 560 190 580
rect 150 550 190 560
rect 105 515 130 530
rect 115 505 130 515
rect 50 350 65 405
rect 115 350 130 405
rect 50 240 65 250
rect 15 225 65 240
rect 15 130 30 225
rect 115 210 130 250
rect 80 195 130 210
rect 55 185 95 195
rect 55 165 65 185
rect 85 165 95 185
rect 55 155 95 165
rect 120 160 160 170
rect 120 140 130 160
rect 150 140 160 160
rect 120 130 160 140
rect 15 115 65 130
rect 50 105 65 115
rect 115 115 135 130
rect 115 105 130 115
rect 50 -10 65 5
rect 115 -10 130 5
rect 25 -20 65 -10
rect 25 -40 35 -20
rect 55 -40 65 -20
rect 25 -50 65 -40
<< polycont >>
rect 30 1650 50 1670
rect 95 1635 115 1655
rect 0 1225 20 1245
rect 65 1205 85 1225
rect 50 945 70 965
rect 110 780 130 800
rect 95 575 115 595
rect 160 560 180 580
rect 65 165 85 185
rect 130 140 150 160
rect 35 -40 55 -20
<< locali >>
rect -65 1815 -20 1825
rect -65 1745 -50 1815
rect -30 1745 -20 1815
rect -65 1735 -20 1745
rect 5 1815 45 1825
rect 5 1745 15 1815
rect 35 1745 45 1815
rect 5 1735 45 1745
rect 70 1815 110 1825
rect 70 1745 80 1815
rect 100 1745 110 1815
rect 70 1735 110 1745
rect 150 1815 190 1825
rect 150 1745 160 1815
rect 180 1745 190 1815
rect 150 1735 190 1745
rect -40 1575 -20 1735
rect 70 1715 90 1735
rect 40 1695 90 1715
rect 40 1680 60 1695
rect 20 1670 60 1680
rect 20 1650 30 1670
rect 50 1650 60 1670
rect 20 1640 60 1650
rect 85 1655 125 1665
rect 85 1635 95 1655
rect 115 1635 125 1655
rect 85 1625 125 1635
rect 90 1575 110 1625
rect -60 1565 -20 1575
rect -60 1495 -50 1565
rect -30 1495 -20 1565
rect -60 1485 -20 1495
rect 5 1565 45 1575
rect 5 1495 15 1565
rect 35 1495 45 1565
rect 5 1485 45 1495
rect 70 1565 110 1575
rect 70 1495 80 1565
rect 100 1495 110 1565
rect 70 1485 110 1495
rect 70 1460 90 1485
rect 25 1440 90 1460
rect 25 1410 45 1440
rect -85 1400 -20 1410
rect -85 1385 -50 1400
rect -60 1330 -50 1385
rect -30 1330 -20 1400
rect -60 1320 -20 1330
rect 5 1400 45 1410
rect 5 1330 15 1400
rect 35 1330 45 1400
rect 5 1320 45 1330
rect 70 1400 110 1410
rect 70 1330 80 1400
rect 100 1330 110 1400
rect 70 1320 110 1330
rect 130 1390 205 1410
rect 25 1295 45 1320
rect 25 1275 75 1295
rect -10 1245 30 1255
rect -10 1225 0 1245
rect 20 1225 30 1245
rect -10 1215 30 1225
rect 10 1160 30 1215
rect 55 1235 75 1275
rect 55 1225 95 1235
rect 55 1205 65 1225
rect 85 1205 95 1225
rect 55 1195 95 1205
rect -85 1150 -20 1160
rect -85 1135 -50 1150
rect -60 1080 -50 1135
rect -30 1080 -20 1150
rect -60 1070 -20 1080
rect 5 1150 45 1160
rect 5 1080 15 1150
rect 35 1080 45 1150
rect 5 1070 45 1080
rect 70 1150 110 1160
rect 70 1080 80 1150
rect 100 1080 110 1150
rect 70 1070 110 1080
rect 5 1015 25 1070
rect 130 1050 150 1390
rect -80 995 25 1015
rect 100 1030 150 1050
rect 170 1140 205 1160
rect -80 140 -60 995
rect 40 965 80 975
rect 40 955 50 965
rect -40 945 50 955
rect 70 945 80 965
rect -40 935 80 945
rect -40 345 -20 935
rect 100 915 120 1030
rect 100 895 125 915
rect 40 870 80 885
rect 40 810 50 870
rect 70 810 80 870
rect 40 795 80 810
rect 100 810 120 895
rect 100 800 140 810
rect 100 780 110 800
rect 130 780 140 800
rect 100 770 140 780
rect 170 750 190 1140
rect 0 740 45 750
rect 0 670 15 740
rect 35 670 45 740
rect 0 660 45 670
rect 70 740 110 750
rect 70 670 80 740
rect 100 670 110 740
rect 70 660 110 670
rect 135 740 190 750
rect 135 670 145 740
rect 165 730 190 740
rect 165 670 175 730
rect 135 660 175 670
rect 25 500 45 660
rect 135 640 155 660
rect 105 620 155 640
rect 105 605 125 620
rect 85 595 125 605
rect 85 575 95 595
rect 115 575 125 595
rect 85 565 125 575
rect 150 580 190 590
rect 150 560 160 580
rect 180 560 190 580
rect 150 550 190 560
rect 155 500 175 550
rect 0 490 45 500
rect 0 420 15 490
rect 35 420 45 490
rect 0 410 45 420
rect 70 490 110 500
rect 70 420 80 490
rect 100 420 110 490
rect 70 410 110 420
rect 135 490 175 500
rect 135 420 145 490
rect 165 420 175 490
rect 135 410 175 420
rect 135 385 155 410
rect 90 365 155 385
rect 90 345 110 365
rect -40 335 45 345
rect -40 325 15 335
rect 5 265 15 325
rect 35 265 45 335
rect 5 255 45 265
rect 70 335 110 345
rect 70 265 80 335
rect 100 265 110 335
rect 70 255 110 265
rect 135 335 175 345
rect 135 265 145 335
rect 165 265 175 335
rect 135 255 175 265
rect 90 235 110 255
rect 90 215 140 235
rect 55 185 95 195
rect 55 165 65 185
rect 85 165 95 185
rect 55 155 95 165
rect -80 120 30 140
rect 10 100 30 120
rect 75 100 95 155
rect 120 170 140 215
rect 120 160 160 170
rect 120 140 130 160
rect 150 140 160 160
rect 120 130 160 140
rect -75 85 -35 100
rect -75 25 -65 85
rect -45 25 -35 85
rect -75 10 -35 25
rect 5 90 45 100
rect 5 20 15 90
rect 35 20 45 90
rect 5 10 45 20
rect 70 90 110 100
rect 70 20 80 90
rect 100 20 110 90
rect 70 10 110 20
rect 135 90 175 100
rect 135 20 145 90
rect 165 20 175 90
rect 135 10 175 20
rect 25 -20 65 -10
rect 25 -30 35 -20
rect -85 -40 35 -30
rect 55 -30 65 -20
rect 55 -40 205 -30
rect -85 -50 205 -40
<< end >>
