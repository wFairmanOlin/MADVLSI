magic
tech sky130A
timestamp 1614264236
<< nwell >>
rect -60 745 265 1330
<< nmos >>
rect 10 545 25 645
rect 50 545 65 645
rect 115 545 130 645
rect 180 545 195 645
rect 10 175 25 275
rect 50 175 65 275
rect 115 175 130 275
rect 180 175 195 275
<< pmos >>
rect 10 1130 25 1230
rect 75 1130 90 1230
rect 140 1130 155 1230
rect 180 1130 195 1230
rect 10 765 25 865
rect 75 765 90 865
rect 140 765 155 865
rect 180 765 195 865
<< ndiff >>
rect -40 630 10 645
rect -40 560 -25 630
rect -5 560 10 630
rect -40 545 10 560
rect 25 545 50 645
rect 65 630 115 645
rect 65 560 80 630
rect 100 560 115 630
rect 65 545 115 560
rect 130 630 180 645
rect 130 560 145 630
rect 165 560 180 630
rect 130 545 180 560
rect 195 630 245 645
rect 195 560 210 630
rect 230 560 245 630
rect 195 545 245 560
rect -40 260 10 275
rect -40 190 -25 260
rect -5 190 10 260
rect -40 175 10 190
rect 25 175 50 275
rect 65 260 115 275
rect 65 190 80 260
rect 100 190 115 260
rect 65 175 115 190
rect 130 260 180 275
rect 130 190 145 260
rect 165 190 180 260
rect 130 175 180 190
rect 195 260 245 275
rect 195 190 210 260
rect 230 190 245 260
rect 195 175 245 190
<< pdiff >>
rect -40 1215 10 1230
rect -40 1145 -25 1215
rect -5 1145 10 1215
rect -40 1130 10 1145
rect 25 1215 75 1230
rect 25 1145 40 1215
rect 60 1145 75 1215
rect 25 1130 75 1145
rect 90 1215 140 1230
rect 90 1145 105 1215
rect 125 1145 140 1215
rect 90 1130 140 1145
rect 155 1130 180 1230
rect 195 1215 245 1230
rect 195 1145 210 1215
rect 230 1145 245 1215
rect 195 1130 245 1145
rect -40 850 10 865
rect -40 780 -25 850
rect -5 780 10 850
rect -40 765 10 780
rect 25 850 75 865
rect 25 780 40 850
rect 60 780 75 850
rect 25 765 75 780
rect 90 850 140 865
rect 90 780 105 850
rect 125 780 140 850
rect 90 765 140 780
rect 155 765 180 865
rect 195 850 245 865
rect 195 780 210 850
rect 230 780 245 850
rect 195 765 245 780
<< ndiffc >>
rect -25 560 -5 630
rect 80 560 100 630
rect 145 560 165 630
rect 210 560 230 630
rect -25 190 -5 260
rect 80 190 100 260
rect 145 190 165 260
rect 210 190 230 260
<< pdiffc >>
rect -25 1145 -5 1215
rect 40 1145 60 1215
rect 105 1145 125 1215
rect 210 1145 230 1215
rect -25 780 -5 850
rect 40 780 60 850
rect 105 780 125 850
rect 210 780 230 850
<< psubdiff >>
rect 55 130 155 145
rect 55 110 70 130
rect 140 110 155 130
rect 55 95 155 110
<< nsubdiff >>
rect 55 1295 155 1310
rect 55 1275 70 1295
rect 140 1275 155 1295
rect 55 1260 155 1275
<< psubdiffcont >>
rect 70 110 140 130
<< nsubdiffcont >>
rect 70 1275 140 1295
<< poly >>
rect 10 1230 25 1245
rect 75 1230 90 1245
rect 140 1230 155 1245
rect 180 1230 195 1245
rect 10 1110 25 1130
rect 75 1110 90 1130
rect 10 1095 30 1110
rect 15 1015 30 1095
rect -5 1000 30 1015
rect 70 1095 90 1110
rect -5 890 10 1000
rect 70 985 85 1095
rect 140 1050 155 1130
rect 180 1080 195 1130
rect 180 1070 225 1080
rect 180 1060 195 1070
rect 45 975 85 985
rect 45 955 55 975
rect 75 955 85 975
rect 45 945 85 955
rect 125 1035 155 1050
rect 185 1050 195 1060
rect 215 1050 225 1070
rect 185 1040 225 1050
rect 125 950 140 1035
rect 165 1000 205 1010
rect 165 980 175 1000
rect 195 980 205 1000
rect 165 970 205 980
rect 125 935 155 950
rect 70 910 110 920
rect 70 890 80 910
rect 100 890 110 910
rect -5 875 25 890
rect 70 880 110 890
rect 10 865 25 875
rect 75 865 90 880
rect 140 865 155 935
rect 190 895 205 970
rect 180 880 205 895
rect 180 865 195 880
rect 10 740 25 765
rect 75 755 90 765
rect -15 730 25 740
rect -15 710 -5 730
rect 15 710 25 730
rect -15 700 25 710
rect 10 645 25 700
rect 50 740 90 755
rect 140 740 155 765
rect 50 645 65 740
rect 115 730 155 740
rect 115 710 125 730
rect 145 710 155 730
rect 115 700 155 710
rect 115 645 130 700
rect 180 645 195 765
rect 10 535 25 545
rect -5 520 25 535
rect -5 365 10 520
rect 50 490 65 545
rect 50 480 90 490
rect 50 460 60 480
rect 80 460 90 480
rect 50 450 90 460
rect 115 430 130 545
rect 35 415 75 425
rect 35 395 45 415
rect 65 395 75 415
rect 35 385 75 395
rect 100 415 130 430
rect -5 350 25 365
rect 10 275 25 350
rect 50 275 65 385
rect 100 335 115 415
rect 180 410 195 545
rect 165 395 195 410
rect 140 385 180 395
rect 140 365 150 385
rect 170 365 180 385
rect 140 355 180 365
rect 100 320 130 335
rect 115 275 130 320
rect 180 320 220 330
rect 180 300 190 320
rect 210 300 220 320
rect 180 290 220 300
rect 180 275 195 290
rect 10 160 25 175
rect 50 160 65 175
rect 115 160 130 175
rect 180 160 195 175
<< polycont >>
rect 55 955 75 975
rect 195 1050 215 1070
rect 175 980 195 1000
rect 80 890 100 910
rect -5 710 15 730
rect 125 710 145 730
rect 60 460 80 480
rect 45 395 65 415
rect 150 365 170 385
rect 190 300 210 320
<< locali >>
rect 60 1295 150 1305
rect 60 1275 70 1295
rect 140 1275 150 1295
rect 60 1265 150 1275
rect -40 1215 5 1225
rect -40 1145 -25 1215
rect -5 1145 5 1215
rect -40 1135 5 1145
rect 30 1215 70 1225
rect 30 1145 40 1215
rect 60 1145 70 1215
rect 30 1135 70 1145
rect 95 1215 135 1225
rect 95 1145 105 1215
rect 125 1145 135 1215
rect 95 1135 135 1145
rect 195 1215 245 1225
rect 195 1145 210 1215
rect 230 1145 245 1215
rect 195 1135 245 1145
rect 50 1025 70 1135
rect 195 1120 215 1135
rect 145 1100 215 1120
rect 50 1005 125 1025
rect 45 975 85 985
rect 45 970 55 975
rect 30 955 55 970
rect 75 955 85 975
rect 30 945 85 955
rect 30 860 50 945
rect 105 920 125 1005
rect 145 1010 165 1100
rect 185 1070 225 1080
rect 185 1050 195 1070
rect 215 1060 225 1070
rect 215 1050 245 1060
rect 185 1040 245 1050
rect 145 1000 205 1010
rect 145 990 175 1000
rect 165 980 175 990
rect 195 980 205 1000
rect 165 970 205 980
rect 70 910 125 920
rect 70 890 80 910
rect 100 900 125 910
rect 100 890 110 900
rect 70 880 110 890
rect 225 860 245 1040
rect -40 850 5 860
rect -40 780 -25 850
rect -5 780 5 850
rect -40 770 5 780
rect 30 850 70 860
rect 30 780 40 850
rect 60 780 70 850
rect 30 770 70 780
rect 95 850 135 860
rect 95 780 105 850
rect 125 780 135 850
rect 95 770 135 780
rect 200 850 245 860
rect 200 780 210 850
rect 230 780 245 850
rect 200 770 245 780
rect -15 730 25 740
rect -15 710 -5 730
rect 15 710 25 730
rect -15 700 25 710
rect 50 675 70 770
rect 115 730 155 740
rect 115 710 125 730
rect 145 710 155 730
rect 115 700 155 710
rect 200 680 220 770
rect 50 655 90 675
rect 70 640 90 655
rect 155 660 220 680
rect 155 640 175 660
rect -35 630 5 640
rect -35 560 -25 630
rect -5 560 5 630
rect -35 550 5 560
rect 70 630 110 640
rect 70 560 80 630
rect 100 560 110 630
rect 70 550 110 560
rect 135 630 175 640
rect 135 560 145 630
rect 165 560 175 630
rect 135 550 175 560
rect 200 630 240 640
rect 200 560 210 630
rect 230 560 240 630
rect 200 550 240 560
rect 70 530 90 550
rect 10 510 90 530
rect 155 530 175 550
rect 155 510 220 530
rect 10 425 30 510
rect 50 480 90 490
rect 50 460 60 480
rect 80 470 90 480
rect 80 460 115 470
rect 50 450 115 460
rect 10 415 75 425
rect 10 405 45 415
rect 35 395 45 405
rect 65 395 75 415
rect 35 385 75 395
rect 95 375 115 450
rect 90 355 115 375
rect 140 385 180 395
rect 140 365 150 385
rect 170 365 180 385
rect 140 355 180 365
rect 90 270 110 355
rect 140 270 160 355
rect 200 330 220 510
rect 180 320 220 330
rect 180 300 190 320
rect 210 300 220 320
rect 180 290 220 300
rect -35 260 5 270
rect -35 190 -25 260
rect -5 190 5 260
rect -35 180 5 190
rect 70 260 110 270
rect 70 190 80 260
rect 100 190 110 260
rect 70 180 110 190
rect 135 260 175 270
rect 135 190 145 260
rect 165 190 175 260
rect 135 180 175 190
rect 200 260 240 270
rect 200 190 210 260
rect 230 190 240 260
rect 200 180 240 190
rect 60 130 150 140
rect 60 110 70 130
rect 140 110 150 130
rect 60 100 150 110
<< viali >>
rect 70 1275 140 1295
rect 105 1145 125 1215
rect 105 780 125 850
rect -5 710 15 730
rect 125 710 145 730
rect -25 560 -5 630
rect 210 560 230 630
rect -25 190 -5 260
rect 210 190 230 260
rect 70 110 140 130
<< metal1 >>
rect -40 1295 245 1310
rect -40 1275 70 1295
rect 140 1275 245 1295
rect -40 1215 245 1275
rect -40 1145 105 1215
rect 125 1145 245 1215
rect -40 850 245 1145
rect -40 780 105 850
rect 125 780 245 850
rect -40 770 245 780
rect -40 730 245 740
rect -40 710 -5 730
rect 15 710 125 730
rect 145 710 245 730
rect -40 675 245 710
rect -40 630 245 645
rect -40 560 -25 630
rect -5 560 210 630
rect 230 560 245 630
rect -40 260 245 560
rect -40 190 -25 260
rect -5 190 210 260
rect 230 190 245 260
rect -40 130 245 190
rect -40 110 70 130
rect 140 110 245 130
rect -40 95 245 110
<< labels >>
rlabel locali 245 815 245 815 3 q
port 3 e
rlabel locali -40 815 -40 815 7 d
port 1 w
rlabel locali 245 1180 245 1180 3 ~q
port 4 e
rlabel locali -40 1180 -40 1180 7 ~d
port 2 w
rlabel metal1 -40 1285 -40 1285 7 vdd
port 6 w
rlabel metal1 -40 705 -40 705 7 phi
port 5 w
rlabel metal1 -40 120 -40 120 7 gnd
port 7 w
<< end >>
