magic
tech sky130A
timestamp 1614110777
<< nwell >>
rect -85 485 215 1440
<< nmos >>
rect 35 1680 50 1780
rect 100 1680 115 1780
rect -15 1475 0 1575
rect 50 1475 65 1575
rect 60 350 75 450
rect 125 350 140 450
rect 10 105 25 205
rect 75 105 90 205
<< pmos >>
rect -15 1310 0 1410
rect 50 1310 65 1410
rect -15 1065 0 1165
rect 50 1065 65 1165
rect 65 755 80 855
rect 130 755 145 855
rect 65 505 80 605
rect 130 505 145 605
<< ndiff >>
rect -15 1765 35 1780
rect -15 1695 0 1765
rect 20 1695 35 1765
rect -15 1680 35 1695
rect 50 1765 100 1780
rect 50 1695 65 1765
rect 85 1695 100 1765
rect 50 1680 100 1695
rect 115 1765 165 1780
rect 115 1695 130 1765
rect 150 1695 165 1765
rect 115 1680 165 1695
rect -65 1560 -15 1575
rect -65 1490 -50 1560
rect -30 1490 -15 1560
rect -65 1475 -15 1490
rect 0 1560 50 1575
rect 0 1490 15 1560
rect 35 1490 50 1560
rect 0 1475 50 1490
rect 65 1560 115 1575
rect 65 1490 80 1560
rect 100 1490 115 1560
rect 65 1475 115 1490
rect 10 435 60 450
rect 10 365 25 435
rect 45 365 60 435
rect 10 350 60 365
rect 75 435 125 450
rect 75 365 90 435
rect 110 365 125 435
rect 75 350 125 365
rect 140 435 190 450
rect 140 365 155 435
rect 175 365 190 435
rect 140 350 190 365
rect -40 190 10 205
rect -40 120 -25 190
rect -5 120 10 190
rect -40 105 10 120
rect 25 190 75 205
rect 25 120 40 190
rect 60 120 75 190
rect 25 105 75 120
rect 90 190 140 205
rect 90 120 105 190
rect 125 120 140 190
rect 90 105 140 120
<< pdiff >>
rect -65 1395 -15 1410
rect -65 1325 -50 1395
rect -30 1325 -15 1395
rect -65 1310 -15 1325
rect 0 1395 50 1410
rect 0 1325 15 1395
rect 35 1325 50 1395
rect 0 1310 50 1325
rect 65 1395 115 1410
rect 65 1325 80 1395
rect 100 1325 115 1395
rect 65 1310 115 1325
rect -65 1150 -15 1165
rect -65 1080 -50 1150
rect -30 1080 -15 1150
rect -65 1065 -15 1080
rect 0 1150 50 1165
rect 0 1080 15 1150
rect 35 1080 50 1150
rect 0 1065 50 1080
rect 65 1150 115 1165
rect 65 1080 80 1150
rect 100 1080 115 1150
rect 65 1065 115 1080
rect 15 840 65 855
rect 15 770 30 840
rect 50 770 65 840
rect 15 755 65 770
rect 80 840 130 855
rect 80 770 95 840
rect 115 770 130 840
rect 80 755 130 770
rect 145 840 195 855
rect 145 770 160 840
rect 180 770 195 840
rect 145 755 195 770
rect 15 590 65 605
rect 15 520 30 590
rect 50 520 65 590
rect 15 505 65 520
rect 80 590 130 605
rect 80 520 95 590
rect 115 520 130 590
rect 80 505 130 520
rect 145 590 195 605
rect 145 520 160 590
rect 180 520 195 590
rect 145 505 195 520
<< ndiffc >>
rect 0 1695 20 1765
rect 65 1695 85 1765
rect 130 1695 150 1765
rect -50 1490 -30 1560
rect 15 1490 35 1560
rect 80 1490 100 1560
rect 25 365 45 435
rect 90 365 110 435
rect 155 365 175 435
rect -25 120 -5 190
rect 40 120 60 190
rect 105 120 125 190
<< pdiffc >>
rect -50 1325 -30 1395
rect 15 1325 35 1395
rect 80 1325 100 1395
rect -50 1080 -30 1150
rect 15 1080 35 1150
rect 80 1080 100 1150
rect 30 770 50 840
rect 95 770 115 840
rect 160 770 180 840
rect 30 520 50 590
rect 95 520 115 590
rect 160 520 180 590
<< psubdiff >>
rect -65 1765 -15 1780
rect -65 1695 -50 1765
rect -30 1695 -15 1765
rect -65 1680 -15 1695
rect 140 190 190 205
rect 140 120 155 190
rect 175 120 190 190
rect 140 105 190 120
<< nsubdiff >>
rect 10 960 110 975
rect 10 940 30 960
rect 90 940 110 960
rect 10 925 110 940
<< psubdiffcont >>
rect -50 1695 -30 1765
rect 155 120 175 190
<< nsubdiffcont >>
rect 30 940 90 960
<< poly >>
rect 35 1780 50 1795
rect 100 1780 115 1795
rect 35 1670 50 1680
rect -15 1655 50 1670
rect -15 1575 0 1655
rect 25 1620 65 1630
rect 100 1625 115 1680
rect 25 1600 35 1620
rect 55 1600 65 1620
rect 25 1590 65 1600
rect 50 1575 65 1590
rect 90 1615 130 1625
rect 90 1595 100 1615
rect 120 1595 130 1615
rect 90 1585 130 1595
rect -15 1410 0 1475
rect 50 1410 65 1475
rect -15 1295 0 1310
rect -50 1280 0 1295
rect -50 1190 -35 1280
rect 50 1260 65 1310
rect 15 1255 65 1260
rect 0 1245 65 1255
rect 0 1225 10 1245
rect 30 1225 40 1245
rect 0 1215 40 1225
rect 65 1210 105 1220
rect 65 1195 75 1210
rect 50 1190 75 1195
rect 95 1190 105 1210
rect -50 1175 0 1190
rect -15 1165 0 1175
rect 50 1180 105 1190
rect 50 1165 65 1180
rect -15 1045 0 1065
rect -60 1030 0 1045
rect 50 1030 65 1065
rect -60 880 -45 1030
rect 50 1020 90 1030
rect 50 1000 60 1020
rect 80 1000 90 1020
rect 50 990 90 1000
rect 110 900 150 910
rect 110 880 120 900
rect 140 880 150 900
rect -60 865 80 880
rect 110 870 150 880
rect 65 855 80 865
rect 130 855 145 870
rect 65 745 80 755
rect 45 730 80 745
rect 130 745 145 755
rect 130 730 170 745
rect 45 630 60 730
rect 85 695 125 705
rect 155 695 170 730
rect 85 675 95 695
rect 115 675 125 695
rect 85 665 125 675
rect 150 685 190 695
rect 150 665 160 685
rect 180 665 190 685
rect 105 630 120 665
rect 150 655 190 665
rect 45 615 80 630
rect 105 615 145 630
rect 65 605 80 615
rect 130 605 145 615
rect 65 495 80 505
rect 130 495 145 505
rect 60 480 80 495
rect 125 480 145 495
rect 60 450 75 480
rect 125 450 140 480
rect 60 340 75 350
rect 10 325 75 340
rect 10 205 25 325
rect 125 300 140 350
rect 50 290 140 300
rect 50 270 60 290
rect 80 285 140 290
rect 80 270 90 285
rect 50 260 90 270
rect 115 250 155 260
rect 115 230 125 250
rect 145 230 155 250
rect 75 220 155 230
rect 75 215 130 220
rect 75 205 90 215
rect 10 90 25 105
rect 75 90 90 105
rect -15 80 25 90
rect -15 60 -5 80
rect 15 60 25 80
rect -15 50 25 60
<< polycont >>
rect 35 1600 55 1620
rect 100 1595 120 1615
rect 10 1225 30 1245
rect 75 1190 95 1210
rect 60 1000 80 1020
rect 120 880 140 900
rect 95 675 115 695
rect 160 665 180 685
rect 60 270 80 290
rect 125 230 145 250
rect -5 60 15 80
<< locali >>
rect -60 1765 30 1775
rect -60 1695 -50 1765
rect -30 1695 0 1765
rect 20 1695 30 1765
rect -60 1685 30 1695
rect 55 1765 95 1775
rect 55 1695 65 1765
rect 85 1695 95 1765
rect 55 1685 95 1695
rect 120 1765 160 1775
rect 120 1695 130 1765
rect 150 1695 160 1765
rect 120 1685 160 1695
rect 120 1665 140 1685
rect 45 1645 140 1665
rect 45 1630 65 1645
rect 25 1620 65 1630
rect 25 1600 35 1620
rect 55 1600 65 1620
rect 25 1590 65 1600
rect 90 1615 130 1625
rect 90 1595 100 1615
rect 120 1595 130 1615
rect 90 1585 130 1595
rect 90 1570 110 1585
rect -60 1560 -20 1570
rect -60 1490 -50 1560
rect -30 1490 -20 1560
rect -60 1480 -20 1490
rect 5 1560 45 1570
rect 5 1490 15 1560
rect 35 1490 45 1560
rect 5 1480 45 1490
rect 70 1560 110 1570
rect 70 1490 80 1560
rect 100 1490 110 1560
rect 70 1480 110 1490
rect 70 1455 90 1480
rect 25 1435 90 1455
rect 25 1405 45 1435
rect -70 1395 -20 1405
rect -70 1385 -50 1395
rect -60 1325 -50 1385
rect -30 1325 -20 1395
rect -60 1315 -20 1325
rect 5 1395 45 1405
rect 5 1325 15 1395
rect 35 1325 45 1395
rect 5 1315 45 1325
rect 70 1395 110 1405
rect 70 1325 80 1395
rect 100 1325 110 1395
rect 70 1315 110 1325
rect 130 1385 205 1405
rect 25 1295 45 1315
rect 25 1275 85 1295
rect 0 1245 40 1255
rect 0 1225 10 1245
rect 30 1225 40 1245
rect 0 1215 40 1225
rect 65 1220 85 1275
rect 10 1160 30 1215
rect 65 1210 105 1220
rect 65 1190 75 1210
rect 95 1190 105 1210
rect 65 1180 105 1190
rect -70 1150 -20 1160
rect -70 1140 -50 1150
rect -60 1080 -50 1140
rect -30 1080 -20 1150
rect -60 1070 -20 1080
rect 5 1150 45 1160
rect 5 1080 15 1150
rect 35 1080 45 1150
rect 5 1070 45 1080
rect 70 1150 110 1160
rect 70 1080 80 1150
rect 100 1080 110 1150
rect 70 1070 110 1080
rect 5 1050 25 1070
rect -65 1030 25 1050
rect -65 200 -45 1030
rect 50 1020 90 1030
rect 50 1010 60 1020
rect -25 1000 60 1010
rect 80 1000 90 1020
rect -25 990 90 1000
rect -25 445 -5 990
rect 15 960 105 970
rect 15 940 30 960
rect 90 940 105 960
rect 15 930 105 940
rect 130 910 150 1385
rect 110 900 150 910
rect 110 880 120 900
rect 140 880 150 900
rect 110 870 150 880
rect 170 1140 205 1160
rect 170 850 190 1140
rect 15 840 60 850
rect 15 770 30 840
rect 50 770 60 840
rect 15 760 60 770
rect 85 840 125 850
rect 85 770 95 840
rect 115 770 125 840
rect 85 760 125 770
rect 150 840 190 850
rect 150 770 160 840
rect 180 770 190 840
rect 150 760 190 770
rect 150 740 170 760
rect 105 720 170 740
rect 105 705 125 720
rect 85 695 125 705
rect 85 675 95 695
rect 115 675 125 695
rect 85 665 125 675
rect 150 685 190 695
rect 150 665 160 685
rect 180 665 190 685
rect 150 655 190 665
rect 160 600 180 655
rect 15 590 60 600
rect 15 520 30 590
rect 50 520 60 590
rect 15 510 60 520
rect 85 590 125 600
rect 85 520 95 590
rect 115 520 125 590
rect 85 510 125 520
rect 150 590 190 600
rect 150 520 160 590
rect 180 520 190 590
rect 150 510 190 520
rect 150 485 170 510
rect 100 465 170 485
rect 100 445 120 465
rect -25 435 55 445
rect -25 425 25 435
rect 15 365 25 425
rect 45 365 55 435
rect 15 355 55 365
rect 80 435 120 445
rect 80 365 90 435
rect 110 365 120 435
rect 80 355 120 365
rect 145 435 185 445
rect 145 365 155 435
rect 175 365 185 435
rect 145 355 185 365
rect 100 335 120 355
rect 100 315 150 335
rect 50 290 90 300
rect 50 270 60 290
rect 80 270 90 290
rect 50 260 90 270
rect 130 260 150 315
rect 50 205 70 260
rect 115 250 155 260
rect 115 230 125 250
rect 145 230 155 250
rect 115 220 155 230
rect 35 200 70 205
rect -65 190 5 200
rect -65 180 -25 190
rect -35 120 -25 180
rect -5 120 5 190
rect -35 110 5 120
rect 30 190 70 200
rect 30 120 40 190
rect 60 120 70 190
rect 30 110 70 120
rect 95 190 185 200
rect 95 120 105 190
rect 125 120 155 190
rect 175 120 185 190
rect 95 110 185 120
rect -15 80 25 90
rect -15 70 -5 80
rect -70 60 -5 70
rect 15 70 25 80
rect 15 60 205 70
rect -70 50 205 60
<< end >>
