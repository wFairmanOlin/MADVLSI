magic
tech sky130A
timestamp 1616204246
<< locali >>
rect 4120 2515 4160 2525
rect 4120 2495 4130 2515
rect 4150 2495 4160 2515
rect 4120 810 4160 2495
rect 4180 1560 4220 1570
rect 4180 1540 4190 1560
rect 4210 1540 4220 1560
rect 4180 865 4220 1540
rect 4180 845 4190 865
rect 4210 845 4220 865
rect 4180 835 4220 845
rect 4120 790 4130 810
rect 4150 790 4160 810
rect 4120 780 4160 790
rect 4070 755 4110 765
rect 4070 735 4080 755
rect 4100 735 4110 755
rect 4070 -10 4110 735
rect 4130 700 4170 710
rect 4130 680 4140 700
rect 4160 680 4170 700
rect 4130 45 4170 680
rect 4130 25 4140 45
rect 4160 25 4170 45
rect 4130 15 4170 25
rect 4070 -30 4080 -10
rect 4100 -30 4110 -10
rect 4070 -40 4110 -30
<< viali >>
rect 4130 2495 4150 2515
rect 4190 1540 4210 1560
rect 4190 845 4210 865
rect 4130 790 4150 810
rect 4080 735 4100 755
rect 4140 680 4160 700
rect 4140 25 4160 45
rect 4080 -30 4100 -10
<< metal1 >>
rect 4120 2515 4220 2525
rect 4120 2495 4130 2515
rect 4150 2495 4220 2515
rect 4120 2485 4220 2495
rect 4180 1560 4220 1570
rect 4180 1540 4190 1560
rect 4210 1540 4220 1560
rect 4180 1530 4220 1540
rect 3895 905 4320 1500
rect 3930 865 4220 875
rect 3930 845 4190 865
rect 4210 845 4220 865
rect 3930 835 4220 845
rect 3960 810 4160 820
rect 3960 790 4130 810
rect 4150 790 4160 810
rect 3960 780 4160 790
rect 3965 755 4110 765
rect 3965 735 4080 755
rect 4100 735 4110 755
rect 3965 725 4110 735
rect 3935 700 4170 710
rect 3935 680 4140 700
rect 4160 680 4170 700
rect 3935 670 4170 680
rect 3875 85 4305 640
rect 4130 45 4225 55
rect 4130 25 4140 45
rect 4160 25 4225 45
rect 4130 15 4225 25
rect 4070 -10 4220 0
rect 4070 -30 4080 -10
rect 4100 -30 4220 -10
rect 4070 -40 4220 -30
use diff_amp  diff_amp_0
timestamp 1616192450
transform 1 0 4445 0 1 -185
box -245 140 1795 2715
use bias_generator  bias_generator_0
timestamp 1616190960
transform 1 0 200 0 1 90
box -220 -100 3770 1470
<< end >>
