magic
tech sky130A
timestamp 1614270699
<< nwell >>
rect -215 275 -50 860
<< nmos >>
rect -145 75 -130 175
<< pmos >>
rect -145 620 -130 720
<< ndiff >>
rect -195 160 -145 175
rect -195 90 -180 160
rect -160 90 -145 160
rect -195 75 -145 90
rect -130 160 -80 175
rect -130 90 -115 160
rect -95 90 -80 160
rect -130 75 -80 90
<< pdiff >>
rect -195 705 -145 720
rect -195 635 -180 705
rect -160 635 -145 705
rect -195 620 -145 635
rect -130 705 -80 720
rect -130 635 -115 705
rect -95 635 -80 705
rect -130 620 -80 635
<< ndiffc >>
rect -180 90 -160 160
rect -115 90 -95 160
<< pdiffc >>
rect -180 635 -160 705
rect -115 635 -95 705
<< psubdiff >>
rect -185 -10 -85 5
rect -185 -30 -170 -10
rect -100 -30 -85 -10
rect -185 -45 -85 -30
<< nsubdiff >>
rect -190 825 -90 840
rect -190 805 -175 825
rect -105 805 -90 825
rect -190 790 -90 805
<< psubdiffcont >>
rect -170 -30 -100 -10
<< nsubdiffcont >>
rect -175 805 -105 825
<< poly >>
rect -145 720 -130 735
rect -145 390 -130 620
rect -145 380 -105 390
rect -145 360 -135 380
rect -115 360 -105 380
rect -145 350 -105 360
rect -145 175 -130 350
rect -145 60 -130 75
rect -170 50 -130 60
rect -170 30 -160 50
rect -140 30 -130 50
rect -170 20 -130 30
<< polycont >>
rect -135 360 -115 380
rect -160 30 -140 50
<< locali >>
rect -185 825 -95 835
rect -185 805 -175 825
rect -105 805 -95 825
rect -185 795 -95 805
rect -170 735 -50 755
rect -170 715 -150 735
rect -195 705 -150 715
rect -195 635 -180 705
rect -160 635 -150 705
rect -195 625 -150 635
rect -125 705 -85 715
rect -125 635 -115 705
rect -95 635 -85 705
rect -125 625 -85 635
rect -185 170 -165 625
rect -145 380 -50 390
rect -145 360 -135 380
rect -115 370 -50 380
rect -115 360 -105 370
rect -145 350 -105 360
rect -190 160 -150 170
rect -190 90 -180 160
rect -160 90 -150 160
rect -190 80 -150 90
rect -125 160 -85 170
rect -125 90 -115 160
rect -95 90 -85 160
rect -125 80 -85 90
rect -215 50 -130 60
rect -215 40 -160 50
rect -170 30 -160 40
rect -140 30 -130 50
rect -170 20 -130 30
rect -180 -10 -90 0
rect -180 -30 -170 -10
rect -100 -30 -90 -10
rect -180 -40 -90 -30
<< viali >>
rect -175 805 -105 825
rect -115 635 -95 705
rect -115 90 -95 160
rect -170 -30 -100 -10
<< metal1 >>
rect -215 825 -50 840
rect -215 805 -175 825
rect -105 805 -50 825
rect -215 705 -50 805
rect -215 635 -115 705
rect -95 635 -50 705
rect -215 300 -50 635
rect -215 205 -50 270
rect -215 160 -50 175
rect -215 90 -115 160
rect -95 90 -50 160
rect -215 -10 -50 90
rect -215 -30 -170 -10
rect -100 -30 -50 -10
rect -215 -55 -50 -30
<< labels >>
rlabel locali -215 50 -215 50 7 d
rlabel metal1 -215 -20 -215 -20 7 gnd
rlabel metal1 -215 240 -215 240 7 phi
rlabel metal1 -215 815 -215 815 7 vdd
rlabel locali -50 745 -50 745 3 ~d
<< end >>
