magic
tech sky130A
timestamp 1612927299
<< nwell >>
rect -380 175 -110 315
<< nmos >>
rect -260 40 -245 140
rect -220 40 -205 140
<< pmos >>
rect -260 195 -245 295
rect -195 195 -180 295
<< ndiff >>
rect -310 130 -260 140
rect -310 50 -295 130
rect -275 50 -260 130
rect -310 40 -260 50
rect -245 40 -220 140
rect -205 130 -155 140
rect -205 50 -190 130
rect -170 50 -155 130
rect -205 40 -155 50
<< pdiff >>
rect -310 285 -260 295
rect -310 205 -295 285
rect -275 205 -260 285
rect -310 195 -260 205
rect -245 285 -195 295
rect -245 205 -230 285
rect -210 205 -195 285
rect -245 195 -195 205
rect -180 285 -130 295
rect -180 205 -165 285
rect -145 205 -130 285
rect -180 195 -130 205
<< ndiffc >>
rect -295 50 -275 130
rect -190 50 -170 130
<< pdiffc >>
rect -295 205 -275 285
rect -230 205 -210 285
rect -165 205 -145 285
<< psubdiff >>
rect -360 130 -310 140
rect -360 50 -345 130
rect -325 50 -310 130
rect -360 40 -310 50
<< nsubdiff >>
rect -360 285 -310 295
rect -360 205 -345 285
rect -325 205 -310 285
rect -360 195 -310 205
<< psubdiffcont >>
rect -345 50 -325 130
<< nsubdiffcont >>
rect -345 205 -325 285
<< poly >>
rect -220 340 -180 350
rect -220 320 -210 340
rect -190 320 -180 340
rect -220 310 -180 320
rect -260 295 -245 310
rect -195 295 -180 310
rect -260 140 -245 195
rect -195 170 -180 195
rect -220 155 -180 170
rect -220 140 -205 155
rect -260 25 -245 40
rect -220 25 -205 40
rect -285 15 -245 25
rect -285 -5 -275 15
rect -255 -5 -245 15
rect -285 -15 -245 -5
<< polycont >>
rect -210 320 -190 340
rect -275 -5 -255 15
<< locali >>
rect -220 340 -180 350
rect -220 330 -210 340
rect -380 320 -210 330
rect -190 320 -180 340
rect -380 310 -180 320
rect -355 285 -265 290
rect -355 205 -345 285
rect -325 205 -295 285
rect -275 205 -265 285
rect -355 200 -265 205
rect -240 285 -200 290
rect -240 205 -230 285
rect -210 205 -200 285
rect -240 200 -200 205
rect -175 285 -130 290
rect -175 205 -165 285
rect -145 205 -130 285
rect -175 200 -130 205
rect -230 175 -210 200
rect -230 155 -165 175
rect -185 135 -165 155
rect -355 130 -265 135
rect -355 50 -345 130
rect -325 50 -295 130
rect -275 50 -265 130
rect -355 45 -265 50
rect -200 130 -160 135
rect -200 50 -190 130
rect -170 50 -160 130
rect -200 45 -160 50
rect -190 25 -170 45
rect -380 15 -245 25
rect -380 5 -275 15
rect -285 -5 -275 5
rect -255 -5 -245 15
rect -190 5 -110 25
rect -285 -15 -245 -5
<< viali >>
rect -345 205 -325 285
rect -295 205 -275 285
rect -165 205 -145 285
rect -345 50 -325 130
rect -295 50 -275 130
<< metal1 >>
rect -380 285 -110 290
rect -380 205 -345 285
rect -325 205 -295 285
rect -275 205 -165 285
rect -145 205 -110 285
rect -380 200 -110 205
rect -380 130 -110 135
rect -380 50 -345 130
rect -325 50 -295 130
rect -275 50 -110 130
rect -380 45 -110 50
<< labels >>
rlabel locali -380 15 -380 15 7 B
port 1 w
rlabel locali -380 320 -380 320 7 A
port 2 w
rlabel metal1 -380 90 -380 90 7 VN
port 4 w
rlabel metal1 -380 245 -380 245 7 VP
port 5 w
rlabel locali -110 15 -110 15 3 Y
port 3 e
<< end >>
