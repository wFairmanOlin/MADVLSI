magic
tech sky130A
timestamp 1616190960
<< nwell >>
rect -220 790 3770 1430
<< nmos >>
rect -100 -45 -50 555
rect 0 -45 50 555
rect 100 -45 150 555
rect 200 -45 250 555
rect 300 -45 350 555
rect 400 -45 450 555
rect 500 -45 550 555
rect 600 -45 650 555
rect 700 -45 750 555
rect 800 -45 850 555
rect 900 -45 950 555
rect 1000 -45 1050 555
rect 1100 -45 1150 555
rect 1200 -45 1250 555
rect 1300 -45 1350 555
rect 1500 -45 1550 555
rect 1600 -45 1650 555
rect 1700 -45 1750 555
rect 1800 -45 1850 555
rect 1900 -45 1950 555
rect 2000 -45 2050 555
rect 2200 -45 2250 555
rect 2300 -45 2350 555
rect 2400 -45 2450 555
rect 2500 -45 2550 555
rect 2600 -45 2650 555
rect 2700 -45 2750 555
rect 2800 -45 2850 555
rect 2900 -45 2950 555
rect 3000 -45 3050 555
rect 3100 -45 3150 555
rect 3200 -45 3250 555
rect 3300 -45 3350 555
rect 3400 -45 3450 555
rect 3500 -45 3550 555
rect 3600 -45 3650 555
<< pmos >>
rect -100 810 -50 1410
rect 0 810 50 1410
rect 100 810 150 1410
rect 200 810 250 1410
rect 300 810 350 1410
rect 400 810 450 1410
rect 500 810 550 1410
rect 600 810 650 1410
rect 700 810 750 1410
rect 800 810 850 1410
rect 900 810 950 1410
rect 1000 810 1050 1410
rect 1100 810 1150 1410
rect 1200 810 1250 1410
rect 1300 810 1350 1410
rect 1500 810 1550 1410
rect 1600 810 1650 1410
rect 1700 810 1750 1410
rect 1800 810 1850 1410
rect 1900 810 1950 1410
rect 2000 810 2050 1410
rect 2200 810 2250 1410
rect 2300 810 2350 1410
rect 2400 810 2450 1410
rect 2500 810 2550 1410
rect 2600 810 2650 1410
rect 2700 810 2750 1410
rect 2800 810 2850 1410
rect 2900 810 2950 1410
rect 3000 810 3050 1410
rect 3100 810 3150 1410
rect 3200 810 3250 1410
rect 3300 810 3350 1410
rect 3400 810 3450 1410
rect 3500 810 3550 1410
rect 3600 810 3650 1410
<< ndiff >>
rect -150 545 -100 555
rect -150 -30 -135 545
rect -115 -30 -100 545
rect -150 -45 -100 -30
rect -50 545 0 555
rect -50 -30 -35 545
rect -15 -30 0 545
rect -50 -45 0 -30
rect 50 545 100 555
rect 50 -30 65 545
rect 85 -30 100 545
rect 50 -45 100 -30
rect 150 545 200 555
rect 150 -30 165 545
rect 185 -30 200 545
rect 150 -45 200 -30
rect 250 545 300 555
rect 250 -30 265 545
rect 285 -30 300 545
rect 250 -45 300 -30
rect 350 545 400 555
rect 350 -30 365 545
rect 385 -30 400 545
rect 350 -45 400 -30
rect 450 545 500 555
rect 450 -30 465 545
rect 485 -30 500 545
rect 450 -45 500 -30
rect 550 545 600 555
rect 550 -30 565 545
rect 585 -30 600 545
rect 550 -45 600 -30
rect 650 545 700 555
rect 650 -30 665 545
rect 685 -30 700 545
rect 650 -45 700 -30
rect 750 545 800 555
rect 750 -30 765 545
rect 785 -30 800 545
rect 750 -45 800 -30
rect 850 545 900 555
rect 850 -30 865 545
rect 885 -30 900 545
rect 850 -45 900 -30
rect 950 545 1000 555
rect 950 -30 965 545
rect 985 -30 1000 545
rect 950 -45 1000 -30
rect 1050 545 1100 555
rect 1050 -30 1065 545
rect 1085 -30 1100 545
rect 1050 -45 1100 -30
rect 1150 545 1200 555
rect 1150 -30 1165 545
rect 1185 -30 1200 545
rect 1150 -45 1200 -30
rect 1250 545 1300 555
rect 1250 -30 1265 545
rect 1285 -30 1300 545
rect 1250 -45 1300 -30
rect 1350 545 1400 555
rect 1450 545 1500 555
rect 1350 -30 1365 545
rect 1385 -30 1400 545
rect 1450 -30 1465 545
rect 1485 -30 1500 545
rect 1350 -45 1400 -30
rect 1450 -45 1500 -30
rect 1550 545 1600 555
rect 1550 -30 1565 545
rect 1585 -30 1600 545
rect 1550 -45 1600 -30
rect 1650 545 1700 555
rect 1650 -30 1665 545
rect 1685 -30 1700 545
rect 1650 -45 1700 -30
rect 1750 545 1800 555
rect 1750 -30 1765 545
rect 1785 -30 1800 545
rect 1750 -45 1800 -30
rect 1850 545 1900 555
rect 1850 -30 1865 545
rect 1885 -30 1900 545
rect 1850 -45 1900 -30
rect 1950 545 2000 555
rect 1950 -30 1965 545
rect 1985 -30 2000 545
rect 1950 -45 2000 -30
rect 2050 545 2100 555
rect 2150 545 2200 555
rect 2050 -30 2065 545
rect 2085 -30 2100 545
rect 2150 -30 2165 545
rect 2185 -30 2200 545
rect 2050 -45 2100 -30
rect 2150 -45 2200 -30
rect 2250 545 2300 555
rect 2250 -30 2265 545
rect 2285 -30 2300 545
rect 2250 -45 2300 -30
rect 2350 545 2400 555
rect 2350 -30 2365 545
rect 2385 -30 2400 545
rect 2350 -45 2400 -30
rect 2450 545 2500 555
rect 2450 -30 2465 545
rect 2485 -30 2500 545
rect 2450 -45 2500 -30
rect 2550 545 2600 555
rect 2550 -30 2565 545
rect 2585 -30 2600 545
rect 2550 -45 2600 -30
rect 2650 545 2700 555
rect 2650 -30 2665 545
rect 2685 -30 2700 545
rect 2650 -45 2700 -30
rect 2750 545 2800 555
rect 2750 -30 2765 545
rect 2785 -30 2800 545
rect 2750 -45 2800 -30
rect 2850 545 2900 555
rect 2850 -30 2865 545
rect 2885 -30 2900 545
rect 2850 -45 2900 -30
rect 2950 545 3000 555
rect 2950 -30 2965 545
rect 2985 -30 3000 545
rect 2950 -45 3000 -30
rect 3050 545 3100 555
rect 3050 -30 3065 545
rect 3085 -30 3100 545
rect 3050 -45 3100 -30
rect 3150 545 3200 555
rect 3150 -30 3165 545
rect 3185 -30 3200 545
rect 3150 -45 3200 -30
rect 3250 545 3300 555
rect 3250 -30 3265 545
rect 3285 -30 3300 545
rect 3250 -45 3300 -30
rect 3350 545 3400 555
rect 3350 -30 3365 545
rect 3385 -30 3400 545
rect 3350 -45 3400 -30
rect 3450 545 3500 555
rect 3450 -30 3465 545
rect 3485 -30 3500 545
rect 3450 -45 3500 -30
rect 3550 545 3600 555
rect 3550 -30 3565 545
rect 3585 -30 3600 545
rect 3550 -45 3600 -30
rect 3650 545 3700 555
rect 3650 -30 3665 545
rect 3685 -30 3700 545
rect 3650 -45 3700 -30
<< pdiff >>
rect -150 1400 -100 1410
rect -150 825 -135 1400
rect -115 825 -100 1400
rect -150 810 -100 825
rect -50 1400 0 1410
rect -50 825 -35 1400
rect -15 825 0 1400
rect -50 810 0 825
rect 50 1400 100 1410
rect 50 825 65 1400
rect 85 825 100 1400
rect 50 810 100 825
rect 150 1400 200 1410
rect 150 825 165 1400
rect 185 825 200 1400
rect 150 810 200 825
rect 250 1400 300 1410
rect 250 825 265 1400
rect 285 825 300 1400
rect 250 810 300 825
rect 350 1400 400 1410
rect 350 825 365 1400
rect 385 825 400 1400
rect 350 810 400 825
rect 450 1400 500 1410
rect 450 825 465 1400
rect 485 825 500 1400
rect 450 810 500 825
rect 550 1400 600 1410
rect 550 825 565 1400
rect 585 825 600 1400
rect 550 810 600 825
rect 650 1400 700 1410
rect 650 825 665 1400
rect 685 825 700 1400
rect 650 810 700 825
rect 750 1400 800 1410
rect 750 825 765 1400
rect 785 825 800 1400
rect 750 810 800 825
rect 850 1400 900 1410
rect 850 825 865 1400
rect 885 825 900 1400
rect 850 810 900 825
rect 950 1400 1000 1410
rect 950 825 965 1400
rect 985 825 1000 1400
rect 950 810 1000 825
rect 1050 1400 1100 1410
rect 1050 825 1065 1400
rect 1085 825 1100 1400
rect 1050 810 1100 825
rect 1150 1400 1200 1410
rect 1150 825 1165 1400
rect 1185 825 1200 1400
rect 1150 810 1200 825
rect 1250 1400 1300 1410
rect 1250 825 1265 1400
rect 1285 825 1300 1400
rect 1250 810 1300 825
rect 1350 1400 1400 1410
rect 1450 1400 1500 1410
rect 1350 825 1365 1400
rect 1385 825 1400 1400
rect 1450 825 1465 1400
rect 1485 825 1500 1400
rect 1350 810 1400 825
rect 1450 810 1500 825
rect 1550 1400 1600 1410
rect 1550 825 1565 1400
rect 1585 825 1600 1400
rect 1550 810 1600 825
rect 1650 1400 1700 1410
rect 1650 825 1665 1400
rect 1685 825 1700 1400
rect 1650 810 1700 825
rect 1750 1400 1800 1410
rect 1750 825 1765 1400
rect 1785 825 1800 1400
rect 1750 810 1800 825
rect 1850 1400 1900 1410
rect 1850 825 1865 1400
rect 1885 825 1900 1400
rect 1850 810 1900 825
rect 1950 1400 2000 1410
rect 1950 825 1965 1400
rect 1985 825 2000 1400
rect 1950 810 2000 825
rect 2050 1400 2100 1410
rect 2150 1400 2200 1410
rect 2050 825 2065 1400
rect 2085 825 2100 1400
rect 2150 825 2165 1400
rect 2185 825 2200 1400
rect 2050 810 2100 825
rect 2150 810 2200 825
rect 2250 1400 2300 1410
rect 2250 825 2265 1400
rect 2285 825 2300 1400
rect 2250 810 2300 825
rect 2350 1400 2400 1410
rect 2350 825 2365 1400
rect 2385 825 2400 1400
rect 2350 810 2400 825
rect 2450 1400 2500 1410
rect 2450 825 2465 1400
rect 2485 825 2500 1400
rect 2450 810 2500 825
rect 2550 1400 2600 1410
rect 2550 825 2565 1400
rect 2585 825 2600 1400
rect 2550 810 2600 825
rect 2650 1400 2700 1410
rect 2650 825 2665 1400
rect 2685 825 2700 1400
rect 2650 810 2700 825
rect 2750 1400 2800 1410
rect 2750 825 2765 1400
rect 2785 825 2800 1400
rect 2750 810 2800 825
rect 2850 1400 2900 1410
rect 2850 825 2865 1400
rect 2885 825 2900 1400
rect 2850 810 2900 825
rect 2950 1400 3000 1410
rect 2950 825 2965 1400
rect 2985 825 3000 1400
rect 2950 810 3000 825
rect 3050 1400 3100 1410
rect 3050 825 3065 1400
rect 3085 825 3100 1400
rect 3050 810 3100 825
rect 3150 1400 3200 1410
rect 3150 825 3165 1400
rect 3185 825 3200 1400
rect 3150 810 3200 825
rect 3250 1400 3300 1410
rect 3250 825 3265 1400
rect 3285 825 3300 1400
rect 3250 810 3300 825
rect 3350 1400 3400 1410
rect 3350 825 3365 1400
rect 3385 825 3400 1400
rect 3350 810 3400 825
rect 3450 1400 3500 1410
rect 3450 825 3465 1400
rect 3485 825 3500 1400
rect 3450 810 3500 825
rect 3550 1400 3600 1410
rect 3550 825 3565 1400
rect 3585 825 3600 1400
rect 3550 810 3600 825
rect 3650 1400 3700 1410
rect 3650 825 3665 1400
rect 3685 825 3700 1400
rect 3650 810 3700 825
<< ndiffc >>
rect -135 -30 -115 545
rect -35 -30 -15 545
rect 65 -30 85 545
rect 165 -30 185 545
rect 265 -30 285 545
rect 365 -30 385 545
rect 465 -30 485 545
rect 565 -30 585 545
rect 665 -30 685 545
rect 765 -30 785 545
rect 865 -30 885 545
rect 965 -30 985 545
rect 1065 -30 1085 545
rect 1165 -30 1185 545
rect 1265 -30 1285 545
rect 1365 -30 1385 545
rect 1465 -30 1485 545
rect 1565 -30 1585 545
rect 1665 -30 1685 545
rect 1765 -30 1785 545
rect 1865 -30 1885 545
rect 1965 -30 1985 545
rect 2065 -30 2085 545
rect 2165 -30 2185 545
rect 2265 -30 2285 545
rect 2365 -30 2385 545
rect 2465 -30 2485 545
rect 2565 -30 2585 545
rect 2665 -30 2685 545
rect 2765 -30 2785 545
rect 2865 -30 2885 545
rect 2965 -30 2985 545
rect 3065 -30 3085 545
rect 3165 -30 3185 545
rect 3265 -30 3285 545
rect 3365 -30 3385 545
rect 3465 -30 3485 545
rect 3565 -30 3585 545
rect 3665 -30 3685 545
<< pdiffc >>
rect -135 825 -115 1400
rect -35 825 -15 1400
rect 65 825 85 1400
rect 165 825 185 1400
rect 265 825 285 1400
rect 365 825 385 1400
rect 465 825 485 1400
rect 565 825 585 1400
rect 665 825 685 1400
rect 765 825 785 1400
rect 865 825 885 1400
rect 965 825 985 1400
rect 1065 825 1085 1400
rect 1165 825 1185 1400
rect 1265 825 1285 1400
rect 1365 825 1385 1400
rect 1465 825 1485 1400
rect 1565 825 1585 1400
rect 1665 825 1685 1400
rect 1765 825 1785 1400
rect 1865 825 1885 1400
rect 1965 825 1985 1400
rect 2065 825 2085 1400
rect 2165 825 2185 1400
rect 2265 825 2285 1400
rect 2365 825 2385 1400
rect 2465 825 2485 1400
rect 2565 825 2585 1400
rect 2665 825 2685 1400
rect 2765 825 2785 1400
rect 2865 825 2885 1400
rect 2965 825 2985 1400
rect 3065 825 3085 1400
rect 3165 825 3185 1400
rect 3265 825 3285 1400
rect 3365 825 3385 1400
rect 3465 825 3485 1400
rect 3565 825 3585 1400
rect 3665 825 3685 1400
<< psubdiff >>
rect -200 545 -150 555
rect -200 -30 -185 545
rect -165 -30 -150 545
rect -200 -45 -150 -30
rect 1400 545 1450 555
rect 1400 -30 1415 545
rect 1435 -30 1450 545
rect 1400 -45 1450 -30
rect 2100 545 2150 555
rect 2100 -30 2115 545
rect 2135 -30 2150 545
rect 2100 -45 2150 -30
rect 3700 545 3750 555
rect 3700 -30 3715 545
rect 3735 -30 3750 545
rect 3700 -45 3750 -30
<< nsubdiff >>
rect -200 1400 -150 1410
rect -200 825 -185 1400
rect -165 825 -150 1400
rect -200 810 -150 825
rect 1400 1400 1450 1410
rect 1400 825 1415 1400
rect 1435 825 1450 1400
rect 1400 810 1450 825
rect 2100 1400 2150 1410
rect 2100 825 2115 1400
rect 2135 825 2150 1400
rect 2100 810 2150 825
rect 3700 1400 3750 1410
rect 3700 825 3715 1400
rect 3735 825 3750 1400
rect 3700 810 3750 825
<< psubdiffcont >>
rect -185 -30 -165 545
rect 1415 -30 1435 545
rect 2115 -30 2135 545
rect 3715 -30 3735 545
<< nsubdiffcont >>
rect -185 825 -165 1400
rect 1415 825 1435 1400
rect 2115 825 2135 1400
rect 3715 825 3735 1400
<< poly >>
rect 600 1455 650 1470
rect 600 1435 615 1455
rect 635 1435 650 1455
rect -100 1410 -50 1430
rect 0 1410 50 1430
rect 100 1410 150 1430
rect 200 1410 250 1430
rect 300 1410 350 1430
rect 400 1410 450 1430
rect 500 1410 550 1430
rect 600 1410 650 1435
rect 1300 1455 1350 1470
rect 1300 1435 1315 1455
rect 1335 1435 1350 1455
rect 700 1410 750 1430
rect 800 1410 850 1430
rect 900 1410 950 1430
rect 1000 1410 1050 1430
rect 1100 1410 1150 1430
rect 1200 1410 1250 1430
rect 1300 1410 1350 1435
rect 1500 1455 1550 1470
rect 1500 1435 1515 1455
rect 1535 1435 1550 1455
rect 1500 1410 1550 1435
rect 1600 1455 1650 1470
rect 1600 1435 1615 1455
rect 1635 1435 1650 1455
rect 1600 1410 1650 1435
rect 1700 1455 1750 1470
rect 1700 1435 1715 1455
rect 1735 1435 1750 1455
rect 1700 1410 1750 1435
rect 1800 1455 1850 1470
rect 1800 1435 1815 1455
rect 1835 1435 1850 1455
rect 1800 1410 1850 1435
rect 1900 1455 1950 1470
rect 1900 1435 1915 1455
rect 1935 1435 1950 1455
rect 1900 1410 1950 1435
rect 2000 1455 2050 1470
rect 2000 1435 2015 1455
rect 2035 1435 2050 1455
rect 2000 1410 2050 1435
rect 2200 1455 2250 1470
rect 2200 1435 2215 1455
rect 2235 1435 2250 1455
rect 2200 1410 2250 1435
rect 2900 1455 2950 1470
rect 2900 1435 2915 1455
rect 2935 1435 2950 1455
rect 2300 1410 2350 1430
rect 2400 1410 2450 1430
rect 2500 1410 2550 1430
rect 2600 1410 2650 1430
rect 2700 1410 2750 1430
rect 2800 1410 2850 1430
rect 2900 1410 2950 1435
rect 3000 1410 3050 1430
rect 3100 1410 3150 1430
rect 3200 1410 3250 1430
rect 3300 1410 3350 1430
rect 3400 1410 3450 1430
rect 3500 1410 3550 1430
rect 3600 1410 3650 1430
rect -100 790 -50 810
rect -150 775 -50 790
rect -150 755 -135 775
rect -115 755 -50 775
rect -150 740 -50 755
rect 0 790 50 810
rect 0 775 60 790
rect 0 755 25 775
rect 45 755 60 775
rect 0 740 60 755
rect 100 775 150 810
rect 100 755 115 775
rect 135 755 150 775
rect 100 740 150 755
rect 200 775 250 810
rect 200 755 215 775
rect 235 755 250 775
rect 200 740 250 755
rect 300 775 350 810
rect 300 755 315 775
rect 335 755 350 775
rect 300 740 350 755
rect 400 775 450 810
rect 500 790 550 810
rect 600 790 650 810
rect 400 755 415 775
rect 435 755 450 775
rect 400 740 450 755
rect 490 775 550 790
rect 490 755 505 775
rect 525 755 550 775
rect 490 740 550 755
rect 700 775 750 810
rect 700 755 715 775
rect 735 755 750 775
rect 700 740 750 755
rect 800 775 850 810
rect 800 755 815 775
rect 835 755 850 775
rect 800 740 850 755
rect 900 775 950 810
rect 900 755 915 775
rect 935 755 950 775
rect 900 740 950 755
rect 1000 775 1050 810
rect 1000 755 1015 775
rect 1035 755 1050 775
rect 1000 740 1050 755
rect 1100 775 1150 810
rect 1100 755 1115 775
rect 1135 755 1150 775
rect 1100 740 1150 755
rect 1200 775 1250 810
rect 1300 790 1350 810
rect 1500 790 1550 810
rect 1600 790 1650 810
rect 1200 755 1215 775
rect 1235 755 1250 775
rect 1200 740 1250 755
rect 1700 775 1750 810
rect 1700 755 1715 775
rect 1735 755 1750 775
rect 1700 740 1750 755
rect 1800 775 1850 810
rect 1900 790 1950 810
rect 2000 790 2050 810
rect 2200 790 2250 810
rect 1800 755 1815 775
rect 1835 755 1850 775
rect 1800 740 1850 755
rect 2300 775 2350 810
rect 2300 755 2315 775
rect 2335 755 2350 775
rect 2300 740 2350 755
rect 2400 775 2450 810
rect 2400 755 2415 775
rect 2435 755 2450 775
rect 2400 740 2450 755
rect 2500 775 2550 810
rect 2500 755 2515 775
rect 2535 755 2550 775
rect 2500 740 2550 755
rect 2600 775 2650 810
rect 2600 755 2615 775
rect 2635 755 2650 775
rect 2600 740 2650 755
rect 2700 775 2750 810
rect 2700 755 2715 775
rect 2735 755 2750 775
rect 2700 740 2750 755
rect 2800 775 2850 810
rect 2900 790 2950 810
rect 3000 790 3050 810
rect 2800 755 2815 775
rect 2835 755 2850 775
rect 2800 740 2850 755
rect 3000 775 3060 790
rect 3000 755 3025 775
rect 3045 755 3060 775
rect 3000 740 3060 755
rect 3100 775 3150 810
rect 3100 755 3115 775
rect 3135 755 3150 775
rect 3100 740 3150 755
rect 3200 775 3250 810
rect 3200 755 3215 775
rect 3235 755 3250 775
rect 3200 740 3250 755
rect 3300 775 3350 810
rect 3300 755 3315 775
rect 3335 755 3350 775
rect 3300 740 3350 755
rect 3400 775 3450 810
rect 3500 790 3550 810
rect 3400 755 3415 775
rect 3435 755 3450 775
rect 3400 740 3450 755
rect 3490 775 3550 790
rect 3490 755 3505 775
rect 3525 755 3550 775
rect 3490 740 3550 755
rect 3600 790 3650 810
rect 3600 775 3700 790
rect 3600 755 3665 775
rect 3685 755 3700 775
rect 3600 740 3700 755
rect 0 605 50 620
rect 0 585 15 605
rect 35 585 50 605
rect -100 555 -50 585
rect 0 555 50 585
rect 100 610 150 625
rect 100 590 115 610
rect 135 590 150 610
rect 100 555 150 590
rect 200 610 250 625
rect 200 590 215 610
rect 235 590 250 610
rect 200 555 250 590
rect 300 610 350 625
rect 300 590 315 610
rect 335 590 350 610
rect 300 555 350 590
rect 400 610 450 625
rect 400 590 415 610
rect 435 590 450 610
rect 400 555 450 590
rect 500 610 550 625
rect 500 590 515 610
rect 535 590 550 610
rect 500 555 550 590
rect 700 610 760 625
rect 700 590 725 610
rect 745 590 760 610
rect 600 555 650 585
rect 700 575 760 590
rect 800 610 850 625
rect 800 590 815 610
rect 835 590 850 610
rect 700 555 750 575
rect 800 555 850 590
rect 900 610 950 625
rect 900 590 915 610
rect 935 590 950 610
rect 900 555 950 590
rect 1000 610 1050 625
rect 1000 590 1015 610
rect 1035 590 1050 610
rect 1000 555 1050 590
rect 1100 610 1150 625
rect 1100 590 1115 610
rect 1135 590 1150 610
rect 1100 555 1150 590
rect 1190 610 1250 625
rect 1190 590 1205 610
rect 1225 590 1250 610
rect 1190 575 1250 590
rect 1600 610 1650 625
rect 1600 590 1615 610
rect 1635 590 1650 610
rect 1200 555 1250 575
rect 1300 555 1350 585
rect 1500 555 1550 585
rect 1600 555 1650 590
rect 1690 610 1750 625
rect 1690 590 1705 610
rect 1725 590 1750 610
rect 1690 575 1750 590
rect 1700 555 1750 575
rect 1800 610 1860 625
rect 1800 590 1825 610
rect 1845 590 1860 610
rect 1800 575 1860 590
rect 1900 610 1950 625
rect 1900 590 1915 610
rect 1935 590 1950 610
rect 1800 555 1850 575
rect 1900 555 1950 590
rect 2300 610 2360 625
rect 2300 590 2325 610
rect 2345 590 2360 610
rect 2000 555 2050 585
rect 2200 555 2250 585
rect 2300 575 2360 590
rect 2400 610 2450 625
rect 2400 590 2415 610
rect 2435 590 2450 610
rect 2300 555 2350 575
rect 2400 555 2450 590
rect 2500 610 2550 625
rect 2500 590 2515 610
rect 2535 590 2550 610
rect 2500 555 2550 590
rect 2600 610 2650 625
rect 2600 590 2615 610
rect 2635 590 2650 610
rect 2600 555 2650 590
rect 2700 610 2750 625
rect 2700 590 2715 610
rect 2735 590 2750 610
rect 2700 555 2750 590
rect 2790 610 2850 625
rect 2790 590 2805 610
rect 2825 590 2850 610
rect 2790 575 2850 590
rect 3000 610 3050 625
rect 3000 590 3015 610
rect 3035 590 3050 610
rect 2800 555 2850 575
rect 2900 555 2950 585
rect 3000 555 3050 590
rect 3100 610 3150 625
rect 3100 590 3115 610
rect 3135 590 3150 610
rect 3100 555 3150 590
rect 3200 610 3250 625
rect 3200 590 3215 610
rect 3235 590 3250 610
rect 3200 555 3250 590
rect 3300 610 3350 625
rect 3300 590 3315 610
rect 3335 590 3350 610
rect 3300 555 3350 590
rect 3400 610 3450 625
rect 3400 590 3415 610
rect 3435 590 3450 610
rect 3400 555 3450 590
rect 3500 605 3550 620
rect 3500 585 3515 605
rect 3535 585 3550 605
rect 3500 555 3550 585
rect 3600 555 3650 585
rect -100 -65 -50 -45
rect 0 -65 50 -45
rect 100 -65 150 -45
rect 200 -65 250 -45
rect 300 -65 350 -45
rect 400 -65 450 -45
rect 500 -65 550 -45
rect 600 -65 650 -45
rect 700 -65 750 -45
rect 800 -65 850 -45
rect 900 -65 950 -45
rect 1000 -65 1050 -45
rect 1100 -65 1150 -45
rect 1200 -65 1250 -45
rect 1300 -65 1350 -45
rect -100 -85 -85 -65
rect -65 -85 -50 -65
rect -100 -100 -50 -85
rect 600 -85 615 -65
rect 635 -85 650 -65
rect 600 -100 650 -85
rect 1300 -85 1315 -65
rect 1335 -85 1350 -65
rect 1300 -100 1350 -85
rect 1500 -65 1550 -45
rect 1600 -65 1650 -45
rect 1700 -65 1750 -45
rect 1800 -65 1850 -45
rect 1900 -65 1950 -45
rect 2000 -65 2050 -45
rect 1500 -85 1515 -65
rect 1535 -85 1550 -65
rect 1500 -100 1550 -85
rect 2000 -85 2015 -65
rect 2035 -85 2050 -65
rect 2000 -100 2050 -85
rect 2200 -65 2250 -45
rect 2300 -65 2350 -45
rect 2400 -65 2450 -45
rect 2500 -65 2550 -45
rect 2600 -65 2650 -45
rect 2700 -65 2750 -45
rect 2800 -65 2850 -45
rect 2900 -65 2950 -45
rect 3000 -65 3050 -45
rect 3100 -65 3150 -45
rect 3200 -65 3250 -45
rect 3300 -65 3350 -45
rect 3400 -65 3450 -45
rect 3500 -65 3550 -45
rect 3600 -65 3650 -45
rect 2200 -85 2215 -65
rect 2235 -85 2250 -65
rect 2200 -100 2250 -85
rect 2900 -85 2915 -65
rect 2935 -85 2950 -65
rect 2900 -100 2950 -85
rect 3600 -85 3615 -65
rect 3635 -85 3650 -65
rect 3600 -100 3650 -85
<< polycont >>
rect 615 1435 635 1455
rect 1315 1435 1335 1455
rect 1515 1435 1535 1455
rect 1615 1435 1635 1455
rect 1715 1435 1735 1455
rect 1815 1435 1835 1455
rect 1915 1435 1935 1455
rect 2015 1435 2035 1455
rect 2215 1435 2235 1455
rect 2915 1435 2935 1455
rect -135 755 -115 775
rect 25 755 45 775
rect 115 755 135 775
rect 215 755 235 775
rect 315 755 335 775
rect 415 755 435 775
rect 505 755 525 775
rect 715 755 735 775
rect 815 755 835 775
rect 915 755 935 775
rect 1015 755 1035 775
rect 1115 755 1135 775
rect 1215 755 1235 775
rect 1715 755 1735 775
rect 1815 755 1835 775
rect 2315 755 2335 775
rect 2415 755 2435 775
rect 2515 755 2535 775
rect 2615 755 2635 775
rect 2715 755 2735 775
rect 2815 755 2835 775
rect 3025 755 3045 775
rect 3115 755 3135 775
rect 3215 755 3235 775
rect 3315 755 3335 775
rect 3415 755 3435 775
rect 3505 755 3525 775
rect 3665 755 3685 775
rect 15 585 35 605
rect 115 590 135 610
rect 215 590 235 610
rect 315 590 335 610
rect 415 590 435 610
rect 515 590 535 610
rect 725 590 745 610
rect 815 590 835 610
rect 915 590 935 610
rect 1015 590 1035 610
rect 1115 590 1135 610
rect 1205 590 1225 610
rect 1615 590 1635 610
rect 1705 590 1725 610
rect 1825 590 1845 610
rect 1915 590 1935 610
rect 2325 590 2345 610
rect 2415 590 2435 610
rect 2515 590 2535 610
rect 2615 590 2635 610
rect 2715 590 2735 610
rect 2805 590 2825 610
rect 3015 590 3035 610
rect 3115 590 3135 610
rect 3215 590 3235 610
rect 3315 590 3335 610
rect 3415 590 3435 610
rect 3515 585 3535 605
rect -85 -85 -65 -65
rect 615 -85 635 -65
rect 1315 -85 1335 -65
rect 1515 -85 1535 -65
rect 2015 -85 2035 -65
rect 2215 -85 2235 -65
rect 2915 -85 2935 -65
rect 3615 -85 3635 -65
<< locali >>
rect 605 1455 695 1465
rect 605 1435 615 1455
rect 635 1435 695 1455
rect 605 1425 695 1435
rect -195 1400 -105 1405
rect -195 825 -185 1400
rect -165 825 -135 1400
rect -115 825 -105 1400
rect -195 815 -105 825
rect -145 775 -105 815
rect -145 755 -135 775
rect -115 755 -105 775
rect -145 745 -105 755
rect -45 1400 -5 1405
rect -45 825 -35 1400
rect -15 825 -5 1400
rect -45 665 -5 825
rect 55 1400 95 1405
rect 55 825 65 1400
rect 85 825 95 1400
rect 55 815 95 825
rect 155 1400 195 1405
rect 155 825 165 1400
rect 185 825 195 1400
rect 155 815 195 825
rect 255 1400 295 1405
rect 255 825 265 1400
rect 285 825 295 1400
rect 255 815 295 825
rect 355 1400 395 1405
rect 355 825 365 1400
rect 385 825 395 1400
rect 355 815 395 825
rect 455 1400 495 1405
rect 455 825 465 1400
rect 485 825 495 1400
rect 455 815 495 825
rect 555 1400 595 1405
rect 555 825 565 1400
rect 585 825 595 1400
rect 15 775 55 785
rect 15 755 25 775
rect 45 755 55 775
rect 15 745 55 755
rect 105 775 145 785
rect 105 755 115 775
rect 135 755 145 775
rect 105 745 145 755
rect 205 775 245 785
rect 205 755 215 775
rect 235 755 245 775
rect 205 745 245 755
rect 305 775 345 785
rect 305 755 315 775
rect 335 755 345 775
rect 305 745 345 755
rect 405 775 445 785
rect 405 755 415 775
rect 435 755 445 775
rect 405 745 445 755
rect 495 775 535 785
rect 495 755 505 775
rect 525 755 535 775
rect 495 745 535 755
rect -45 645 -35 665
rect -15 645 -5 665
rect -45 615 -5 645
rect 555 620 595 825
rect 655 1400 695 1425
rect 655 825 665 1400
rect 685 825 695 1400
rect 655 815 695 825
rect 755 1425 1195 1465
rect 1305 1455 1645 1465
rect 1305 1435 1315 1455
rect 1335 1435 1515 1455
rect 1535 1435 1615 1455
rect 1635 1435 1645 1455
rect 1305 1425 1645 1435
rect 1705 1455 1845 1465
rect 1705 1435 1715 1455
rect 1735 1435 1815 1455
rect 1835 1435 1845 1455
rect 1705 1425 1845 1435
rect 1905 1455 2245 1465
rect 1905 1435 1915 1455
rect 1935 1435 2015 1455
rect 2035 1435 2215 1455
rect 2235 1435 2245 1455
rect 1905 1425 2245 1435
rect 2355 1425 2795 1465
rect 755 1400 795 1425
rect 755 825 765 1400
rect 785 825 795 1400
rect 755 815 795 825
rect 855 1400 895 1405
rect 855 825 865 1400
rect 885 825 895 1400
rect 855 785 895 825
rect 955 1400 995 1425
rect 955 825 965 1400
rect 985 825 995 1400
rect 955 815 995 825
rect 1055 1400 1095 1405
rect 1055 825 1065 1400
rect 1085 825 1095 1400
rect 1055 785 1095 825
rect 1155 1400 1195 1425
rect 1155 825 1165 1400
rect 1185 825 1195 1400
rect 1155 815 1195 825
rect 1255 1400 1295 1405
rect 1255 825 1265 1400
rect 1285 825 1295 1400
rect 1255 785 1295 825
rect 1355 1400 1495 1425
rect 1355 825 1365 1400
rect 1385 825 1415 1400
rect 1435 825 1465 1400
rect 1485 825 1495 1400
rect 1355 815 1495 825
rect 1555 1400 1595 1425
rect 1555 825 1565 1400
rect 1585 825 1595 1400
rect 1555 815 1595 825
rect 1655 1400 1695 1410
rect 1655 825 1665 1400
rect 1685 825 1695 1400
rect 1655 815 1695 825
rect 1755 1400 1795 1425
rect 1755 825 1765 1400
rect 1785 825 1795 1400
rect 1755 785 1795 825
rect 1855 1400 1895 1410
rect 1855 825 1865 1400
rect 1885 825 1895 1400
rect 1855 815 1895 825
rect 1955 1400 1995 1425
rect 1955 825 1965 1400
rect 1985 825 1995 1400
rect 1955 815 1995 825
rect 2055 1400 2195 1425
rect 2055 825 2065 1400
rect 2085 825 2115 1400
rect 2135 825 2165 1400
rect 2185 825 2195 1400
rect 2055 815 2195 825
rect 2255 1400 2295 1405
rect 2255 825 2265 1400
rect 2285 825 2295 1400
rect 2255 785 2295 825
rect 2355 1400 2395 1425
rect 2355 825 2365 1400
rect 2385 825 2395 1400
rect 2355 815 2395 825
rect 2455 1400 2495 1405
rect 2455 825 2465 1400
rect 2485 825 2495 1400
rect 2455 785 2495 825
rect 2555 1400 2595 1425
rect 2555 825 2565 1400
rect 2585 825 2595 1400
rect 2555 815 2595 825
rect 2655 1400 2695 1405
rect 2655 825 2665 1400
rect 2685 825 2695 1400
rect 2655 785 2695 825
rect 2755 1400 2795 1425
rect 2755 825 2765 1400
rect 2785 825 2795 1400
rect 2755 815 2795 825
rect 2855 1455 2945 1465
rect 2855 1435 2915 1455
rect 2935 1435 2945 1455
rect 2855 1425 2945 1435
rect 2855 1400 2895 1425
rect 2855 825 2865 1400
rect 2885 825 2895 1400
rect 2855 815 2895 825
rect 2955 1400 2995 1405
rect 2955 825 2965 1400
rect 2985 825 2995 1400
rect -45 605 45 615
rect -45 585 15 605
rect 35 585 45 605
rect -45 575 45 585
rect 105 610 595 620
rect 105 590 115 610
rect 135 590 215 610
rect 235 590 315 610
rect 335 590 415 610
rect 435 590 515 610
rect 535 590 595 610
rect 105 580 595 590
rect 655 775 1145 785
rect 655 755 715 775
rect 735 755 815 775
rect 835 755 915 775
rect 935 755 1015 775
rect 1035 755 1115 775
rect 1135 755 1145 775
rect 655 745 1145 755
rect 1205 775 1295 785
rect 1205 755 1215 775
rect 1235 755 1295 775
rect 1205 745 1295 755
rect 1705 775 1845 785
rect 1705 755 1715 775
rect 1735 755 1815 775
rect 1835 755 1845 775
rect 1705 745 1845 755
rect 2255 775 2345 785
rect 2255 755 2315 775
rect 2335 755 2345 775
rect 2255 745 2345 755
rect 2405 775 2895 785
rect 2405 755 2415 775
rect 2435 755 2515 775
rect 2535 755 2615 775
rect 2635 755 2715 775
rect 2735 755 2815 775
rect 2835 755 2895 775
rect 2405 745 2895 755
rect -195 545 -105 550
rect -195 -30 -185 545
rect -165 -30 -135 545
rect -115 -30 -105 545
rect -195 -40 -105 -30
rect -45 545 -5 575
rect -45 -30 -35 545
rect -15 -30 -5 545
rect -45 -40 -5 -30
rect 55 545 95 550
rect 55 -30 65 545
rect 85 -30 95 545
rect -150 -55 -105 -40
rect -150 -65 -55 -55
rect -150 -85 -85 -65
rect -65 -85 -55 -65
rect -150 -95 -55 -85
rect 55 -60 95 -30
rect 155 545 195 580
rect 155 -30 165 545
rect 185 -30 195 545
rect 155 -40 195 -30
rect 255 545 295 550
rect 255 -30 265 545
rect 285 -30 295 545
rect 255 -60 295 -30
rect 355 545 395 580
rect 355 -30 365 545
rect 385 -30 395 545
rect 355 -40 395 -30
rect 455 545 495 550
rect 455 -30 465 545
rect 485 -30 495 545
rect 455 -60 495 -30
rect 55 -100 495 -60
rect 555 545 595 550
rect 555 -30 565 545
rect 585 -30 595 545
rect 555 -55 595 -30
rect 655 545 695 745
rect 1255 720 1295 745
rect 1255 700 1265 720
rect 1285 700 1295 720
rect 715 610 755 620
rect 715 590 725 610
rect 745 590 755 610
rect 715 580 755 590
rect 805 610 845 620
rect 805 590 815 610
rect 835 590 845 610
rect 805 580 845 590
rect 905 610 945 620
rect 905 590 915 610
rect 935 590 945 610
rect 905 580 945 590
rect 1005 610 1045 620
rect 1005 590 1015 610
rect 1035 590 1045 610
rect 1005 580 1045 590
rect 1105 610 1145 620
rect 1105 590 1115 610
rect 1135 590 1145 610
rect 1105 580 1145 590
rect 1195 610 1235 620
rect 1195 590 1205 610
rect 1225 590 1235 610
rect 1195 580 1235 590
rect 655 -30 665 545
rect 685 -30 695 545
rect 655 -40 695 -30
rect 755 545 795 550
rect 755 -30 765 545
rect 785 -30 795 545
rect 755 -40 795 -30
rect 855 545 895 550
rect 855 -30 865 545
rect 885 -30 895 545
rect 855 -40 895 -30
rect 955 545 995 550
rect 955 -30 965 545
rect 985 -30 995 545
rect 955 -40 995 -30
rect 1055 545 1095 550
rect 1055 -30 1065 545
rect 1085 -30 1095 545
rect 1055 -40 1095 -30
rect 1155 545 1195 550
rect 1155 -30 1165 545
rect 1185 -30 1195 545
rect 1155 -40 1195 -30
rect 1255 545 1295 700
rect 1555 610 1645 620
rect 1555 590 1565 610
rect 1585 590 1615 610
rect 1635 590 1645 610
rect 1555 580 1645 590
rect 1695 610 1735 620
rect 1695 590 1705 610
rect 1725 590 1735 610
rect 1695 580 1735 590
rect 1255 -30 1265 545
rect 1285 -30 1295 545
rect 1255 -40 1295 -30
rect 1355 545 1495 550
rect 1355 -30 1365 545
rect 1385 -30 1415 545
rect 1435 -30 1465 545
rect 1485 -30 1495 545
rect 1355 -55 1495 -30
rect 1555 545 1595 580
rect 1555 -30 1565 545
rect 1585 -30 1595 545
rect 1555 -40 1595 -30
rect 1655 545 1695 550
rect 1655 -30 1665 545
rect 1685 -30 1695 545
rect 1655 -40 1695 -30
rect 1755 545 1795 745
rect 2255 720 2295 745
rect 2255 700 2265 720
rect 2285 700 2295 720
rect 1815 610 1855 620
rect 1815 590 1825 610
rect 1845 590 1855 610
rect 1815 580 1855 590
rect 1905 610 1995 620
rect 1905 590 1915 610
rect 1935 590 1965 610
rect 1985 590 1995 610
rect 1905 580 1995 590
rect 1755 -30 1765 545
rect 1785 -30 1795 545
rect 1755 -40 1795 -30
rect 1855 545 1895 550
rect 1855 -30 1865 545
rect 1885 -30 1895 545
rect 1855 -40 1895 -30
rect 1955 545 1995 580
rect 1955 -30 1965 545
rect 1985 -30 1995 545
rect 1955 -40 1995 -30
rect 2055 545 2195 550
rect 2055 -30 2065 545
rect 2085 -30 2115 545
rect 2135 -30 2165 545
rect 2185 -30 2195 545
rect 2055 -55 2195 -30
rect 2255 545 2295 700
rect 2315 610 2355 620
rect 2315 590 2325 610
rect 2345 590 2355 610
rect 2315 580 2355 590
rect 2405 610 2445 620
rect 2405 590 2415 610
rect 2435 590 2445 610
rect 2405 580 2445 590
rect 2505 610 2545 620
rect 2505 590 2515 610
rect 2535 590 2545 610
rect 2505 580 2545 590
rect 2605 610 2645 620
rect 2605 590 2615 610
rect 2635 590 2645 610
rect 2605 580 2645 590
rect 2705 610 2745 620
rect 2705 590 2715 610
rect 2735 590 2745 610
rect 2705 580 2745 590
rect 2795 610 2835 620
rect 2795 590 2805 610
rect 2825 590 2835 610
rect 2795 580 2835 590
rect 2255 -30 2265 545
rect 2285 -30 2295 545
rect 2255 -40 2295 -30
rect 2355 545 2395 550
rect 2355 -30 2365 545
rect 2385 -30 2395 545
rect 2355 -40 2395 -30
rect 2455 545 2495 550
rect 2455 -30 2465 545
rect 2485 -30 2495 545
rect 2455 -40 2495 -30
rect 2555 545 2595 550
rect 2555 -30 2565 545
rect 2585 -30 2595 545
rect 2555 -40 2595 -30
rect 2655 545 2695 550
rect 2655 -30 2665 545
rect 2685 -30 2695 545
rect 2655 -40 2695 -30
rect 2755 545 2795 550
rect 2755 -30 2765 545
rect 2785 -30 2795 545
rect 2755 -40 2795 -30
rect 2855 545 2895 745
rect 2955 620 2995 825
rect 3055 1400 3095 1405
rect 3055 825 3065 1400
rect 3085 825 3095 1400
rect 3055 815 3095 825
rect 3155 1400 3195 1405
rect 3155 825 3165 1400
rect 3185 825 3195 1400
rect 3155 815 3195 825
rect 3255 1400 3295 1405
rect 3255 825 3265 1400
rect 3285 825 3295 1400
rect 3255 815 3295 825
rect 3355 1400 3395 1405
rect 3355 825 3365 1400
rect 3385 825 3395 1400
rect 3355 815 3395 825
rect 3455 1400 3495 1405
rect 3455 825 3465 1400
rect 3485 825 3495 1400
rect 3455 815 3495 825
rect 3555 1400 3595 1405
rect 3555 825 3565 1400
rect 3585 825 3595 1400
rect 3015 775 3055 785
rect 3015 755 3025 775
rect 3045 755 3055 775
rect 3015 745 3055 755
rect 3105 775 3145 785
rect 3105 755 3115 775
rect 3135 755 3145 775
rect 3105 745 3145 755
rect 3205 775 3245 785
rect 3205 755 3215 775
rect 3235 755 3245 775
rect 3205 745 3245 755
rect 3305 775 3345 785
rect 3305 755 3315 775
rect 3335 755 3345 775
rect 3305 745 3345 755
rect 3405 775 3445 785
rect 3405 755 3415 775
rect 3435 755 3445 775
rect 3405 745 3445 755
rect 3495 775 3535 785
rect 3495 755 3505 775
rect 3525 755 3535 775
rect 3495 745 3535 755
rect 3555 665 3595 825
rect 3655 1400 3745 1405
rect 3655 825 3665 1400
rect 3685 825 3715 1400
rect 3735 825 3745 1400
rect 3655 815 3745 825
rect 3655 775 3695 815
rect 3655 755 3665 775
rect 3685 755 3695 775
rect 3655 745 3695 755
rect 3555 645 3565 665
rect 3585 645 3595 665
rect 2955 610 3445 620
rect 3555 615 3595 645
rect 2955 590 3015 610
rect 3035 590 3115 610
rect 3135 590 3215 610
rect 3235 590 3315 610
rect 3335 590 3415 610
rect 3435 590 3445 610
rect 2955 580 3445 590
rect 3505 605 3595 615
rect 3505 585 3515 605
rect 3535 585 3595 605
rect 2855 -30 2865 545
rect 2885 -30 2895 545
rect 2855 -40 2895 -30
rect 2955 545 2995 550
rect 2955 -30 2965 545
rect 2985 -30 2995 545
rect 2955 -55 2995 -30
rect 555 -65 645 -55
rect 555 -85 615 -65
rect 635 -85 645 -65
rect 555 -95 645 -85
rect 1305 -65 1545 -55
rect 1305 -85 1315 -65
rect 1335 -85 1515 -65
rect 1535 -85 1545 -65
rect 1305 -95 1545 -85
rect 2005 -65 2245 -55
rect 2005 -85 2015 -65
rect 2035 -85 2215 -65
rect 2235 -85 2245 -65
rect 2005 -95 2245 -85
rect 2905 -65 2995 -55
rect 2905 -85 2915 -65
rect 2935 -85 2995 -65
rect 2905 -95 2995 -85
rect 3055 545 3095 550
rect 3055 -30 3065 545
rect 3085 -30 3095 545
rect 3055 -60 3095 -30
rect 3155 545 3195 580
rect 3155 -30 3165 545
rect 3185 -30 3195 545
rect 3155 -40 3195 -30
rect 3255 545 3295 550
rect 3255 -30 3265 545
rect 3285 -30 3295 545
rect 3255 -60 3295 -30
rect 3355 545 3395 580
rect 3505 575 3595 585
rect 3355 -30 3365 545
rect 3385 -30 3395 545
rect 3355 -40 3395 -30
rect 3455 545 3495 550
rect 3455 -30 3465 545
rect 3485 -30 3495 545
rect 3455 -60 3495 -30
rect 3555 545 3595 575
rect 3555 -30 3565 545
rect 3585 -30 3595 545
rect 3555 -40 3595 -30
rect 3655 545 3745 550
rect 3655 -30 3665 545
rect 3685 -30 3715 545
rect 3735 -30 3745 545
rect 3655 -40 3745 -30
rect 3655 -55 3700 -40
rect 3055 -100 3495 -60
rect 3605 -65 3700 -55
rect 3605 -85 3615 -65
rect 3635 -85 3700 -65
rect 3605 -95 3700 -85
<< viali >>
rect -185 825 -165 1400
rect -135 825 -115 1400
rect 65 825 85 1400
rect 25 755 45 775
rect 115 755 135 775
rect 215 755 235 775
rect 315 755 335 775
rect 415 755 435 775
rect 505 755 525 775
rect -35 645 -15 665
rect 665 825 685 1400
rect 1365 825 1385 1400
rect 1415 825 1435 1400
rect 1465 825 1485 1400
rect 1565 825 1585 1400
rect 1665 825 1685 1400
rect 1865 825 1885 1400
rect 1965 825 1985 1400
rect 2065 825 2085 1400
rect 2115 825 2135 1400
rect 2165 825 2185 1400
rect 2865 825 2885 1400
rect 1715 755 1735 775
rect 1815 755 1835 775
rect -185 -30 -165 545
rect -135 -30 -115 545
rect 565 -30 585 545
rect 1265 700 1285 720
rect 725 590 745 610
rect 815 590 835 610
rect 915 590 935 610
rect 1015 590 1035 610
rect 1115 590 1135 610
rect 1205 590 1225 610
rect 1165 -30 1185 545
rect 1565 590 1585 610
rect 1615 590 1635 610
rect 1705 590 1725 610
rect 1365 -30 1385 545
rect 1415 -30 1435 545
rect 1465 -30 1485 545
rect 1665 -30 1685 545
rect 2265 700 2285 720
rect 1825 590 1845 610
rect 1915 590 1935 610
rect 1965 590 1985 610
rect 1865 -30 1885 545
rect 2065 -30 2085 545
rect 2115 -30 2135 545
rect 2165 -30 2185 545
rect 2325 590 2345 610
rect 2415 590 2435 610
rect 2515 590 2535 610
rect 2615 590 2635 610
rect 2715 590 2735 610
rect 2805 590 2825 610
rect 2365 -30 2385 545
rect 3465 825 3485 1400
rect 3025 755 3045 775
rect 3115 755 3135 775
rect 3215 755 3235 775
rect 3315 755 3335 775
rect 3415 755 3435 775
rect 3505 755 3525 775
rect 3665 825 3685 1400
rect 3715 825 3735 1400
rect 3565 645 3585 665
rect 2965 -30 2985 545
rect 3665 -30 3685 545
rect 3715 -30 3735 545
<< metal1 >>
rect -220 1400 3770 1410
rect -220 825 -185 1400
rect -165 825 -135 1400
rect -115 825 65 1400
rect 85 825 665 1400
rect 685 825 1365 1400
rect 1385 825 1415 1400
rect 1435 825 1465 1400
rect 1485 825 1565 1400
rect 1585 825 1665 1400
rect 1685 825 1865 1400
rect 1885 825 1965 1400
rect 1985 825 2065 1400
rect 2085 825 2115 1400
rect 2135 825 2165 1400
rect 2185 825 2865 1400
rect 2885 825 3465 1400
rect 3485 825 3665 1400
rect 3685 825 3715 1400
rect 3735 825 3770 1400
rect -220 815 3770 825
rect -220 775 3770 785
rect -220 755 25 775
rect 45 755 115 775
rect 135 755 215 775
rect 235 755 315 775
rect 335 755 415 775
rect 435 755 505 775
rect 525 755 1715 775
rect 1735 755 1815 775
rect 1835 755 3025 775
rect 3045 755 3115 775
rect 3135 755 3215 775
rect 3235 755 3315 775
rect 3335 755 3415 775
rect 3435 755 3505 775
rect 3525 755 3770 775
rect -220 745 3770 755
rect -220 720 3770 730
rect -220 700 1265 720
rect 1285 700 2265 720
rect 2285 700 3770 720
rect -220 690 3770 700
rect -220 665 3770 675
rect -220 645 -35 665
rect -15 645 3565 665
rect 3585 645 3770 665
rect -220 635 3770 645
rect -220 610 3770 620
rect -220 590 725 610
rect 745 590 815 610
rect 835 590 915 610
rect 935 590 1015 610
rect 1035 590 1115 610
rect 1135 590 1205 610
rect 1225 590 1565 610
rect 1585 590 1615 610
rect 1635 590 1705 610
rect 1725 590 1825 610
rect 1845 590 1915 610
rect 1935 590 1965 610
rect 1985 590 2325 610
rect 2345 590 2415 610
rect 2435 590 2515 610
rect 2535 590 2615 610
rect 2635 590 2715 610
rect 2735 590 2805 610
rect 2825 590 3770 610
rect -220 580 3770 590
rect -220 545 3770 550
rect -220 -30 -185 545
rect -165 -30 -135 545
rect -115 -30 565 545
rect 585 -30 1165 545
rect 1185 -30 1365 545
rect 1385 -30 1415 545
rect 1435 -30 1465 545
rect 1485 -30 1665 545
rect 1685 -30 1865 545
rect 1885 -30 2065 545
rect 2085 -30 2115 545
rect 2135 -30 2165 545
rect 2185 -30 2365 545
rect 2385 -30 2965 545
rect 2985 -30 3665 545
rect 3685 -30 3715 545
rect 3735 -30 3770 545
rect -220 -40 3770 -30
<< labels >>
rlabel metal1 -220 815 -200 1410 7 VDD
rlabel metal1 -220 745 -180 785 7 vbp
rlabel metal1 -220 690 -180 730 7 vcp
rlabel metal1 -220 635 -180 675 7 vcn
rlabel metal1 -220 580 -180 620 7 vbn
rlabel metal1 -220 -40 -200 550 7 GND
rlabel metal1 3750 815 3770 1410 3 VDD
rlabel metal1 3730 745 3770 785 3 vbp
rlabel metal1 3730 690 3770 730 3 vcp
rlabel metal1 3730 635 3770 675 3 vcn
rlabel metal1 3730 580 3770 620 3 vbn
rlabel metal1 3750 -40 3770 550 3 GND
rlabel locali 165 825 185 1400 1 net13
rlabel locali 265 825 285 1400 1 net14
rlabel locali 365 825 385 1400 1 net15
rlabel locali 465 825 485 1400 1 net24
rlabel locali 565 825 585 1400 1 net17
rlabel locali 765 825 785 1400 1 net1
rlabel locali 865 825 885 1400 1 net2
rlabel locali 765 -30 785 545 1 net6
rlabel locali 865 -30 885 545 1 net5
rlabel locali 965 -30 985 545 1 net4
rlabel locali 1065 -30 1085 545 1 net3
<< end >>
