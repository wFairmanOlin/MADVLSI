magic
tech sky130A
timestamp 1616192450
<< nwell >>
rect -145 2620 -50 2660
rect 1600 2620 1695 2660
rect -235 2150 1785 2620
rect -240 1920 1790 2150
rect -245 1715 1790 1920
rect -240 1070 1790 1715
rect -240 1065 -60 1070
rect 1610 1065 1790 1070
<< nmos >>
rect -100 265 -50 865
rect 0 265 50 865
rect 100 265 150 865
rect 200 265 250 865
rect 400 265 450 865
rect 500 265 550 865
rect 600 265 650 865
rect 700 265 750 865
rect 800 265 850 865
rect 900 265 950 865
rect 1000 265 1050 865
rect 1100 265 1150 865
rect 1300 265 1350 865
rect 1400 265 1450 865
rect 1500 265 1550 865
rect 1600 265 1650 865
<< pmos >>
rect -100 2000 -50 2600
rect 0 2000 50 2600
rect 100 2000 150 2600
rect 200 2000 250 2600
rect 400 2000 450 2600
rect 500 2000 550 2600
rect 600 2000 650 2600
rect 700 2000 750 2600
rect 800 2000 850 2600
rect 900 2000 950 2600
rect 1000 2000 1050 2600
rect 1100 2000 1150 2600
rect 1300 2000 1350 2600
rect 1400 2000 1450 2600
rect 1500 2000 1550 2600
rect 1600 2000 1650 2600
rect -95 1090 -45 1690
rect 0 1090 50 1690
rect 100 1090 150 1690
rect 200 1090 250 1690
rect 400 1090 450 1690
rect 500 1090 550 1690
rect 600 1090 650 1690
rect 700 1090 750 1690
rect 800 1090 850 1690
rect 900 1090 950 1690
rect 1000 1090 1050 1690
rect 1100 1090 1150 1690
rect 1300 1090 1350 1690
rect 1400 1090 1450 1690
rect 1500 1090 1550 1690
rect 1595 1090 1645 1690
<< ndiff >>
rect -150 850 -100 865
rect -150 280 -135 850
rect -115 280 -100 850
rect -150 265 -100 280
rect -50 850 0 865
rect -50 280 -35 850
rect -15 280 0 850
rect -50 265 0 280
rect 50 850 100 865
rect 50 280 65 850
rect 85 280 100 850
rect 50 265 100 280
rect 150 850 200 865
rect 150 280 165 850
rect 185 280 200 850
rect 150 265 200 280
rect 250 850 300 865
rect 350 850 400 865
rect 250 280 265 850
rect 285 280 300 850
rect 350 280 365 850
rect 385 280 400 850
rect 250 265 300 280
rect 350 265 400 280
rect 450 850 500 865
rect 450 280 465 850
rect 485 280 500 850
rect 450 265 500 280
rect 550 850 600 865
rect 550 280 565 850
rect 585 280 600 850
rect 550 265 600 280
rect 650 850 700 865
rect 650 280 665 850
rect 685 280 700 850
rect 650 265 700 280
rect 750 850 800 865
rect 750 280 765 850
rect 785 280 800 850
rect 750 265 800 280
rect 850 850 900 865
rect 850 280 865 850
rect 885 280 900 850
rect 850 265 900 280
rect 950 850 1000 865
rect 950 280 965 850
rect 985 280 1000 850
rect 950 265 1000 280
rect 1050 850 1100 865
rect 1050 280 1065 850
rect 1085 280 1100 850
rect 1050 265 1100 280
rect 1150 850 1200 865
rect 1250 850 1300 865
rect 1150 280 1165 850
rect 1185 280 1200 850
rect 1250 280 1265 850
rect 1285 280 1300 850
rect 1150 265 1200 280
rect 1250 265 1300 280
rect 1350 850 1400 865
rect 1350 280 1365 850
rect 1385 280 1400 850
rect 1350 265 1400 280
rect 1450 850 1500 865
rect 1450 280 1465 850
rect 1485 280 1500 850
rect 1450 265 1500 280
rect 1550 850 1600 865
rect 1550 280 1565 850
rect 1585 280 1600 850
rect 1550 265 1600 280
rect 1650 850 1700 865
rect 1650 280 1665 850
rect 1685 280 1700 850
rect 1650 265 1700 280
<< pdiff >>
rect -150 2585 -100 2600
rect -150 2015 -135 2585
rect -115 2015 -100 2585
rect -150 2000 -100 2015
rect -50 2585 0 2600
rect -50 2015 -35 2585
rect -15 2015 0 2585
rect -50 2000 0 2015
rect 50 2585 100 2600
rect 50 2015 65 2585
rect 85 2015 100 2585
rect 50 2000 100 2015
rect 150 2585 200 2600
rect 150 2015 165 2585
rect 185 2015 200 2585
rect 150 2000 200 2015
rect 250 2585 300 2600
rect 350 2585 400 2600
rect 250 2015 265 2585
rect 285 2015 300 2585
rect 350 2015 365 2585
rect 385 2015 400 2585
rect 250 2000 300 2015
rect 350 2000 400 2015
rect 450 2585 500 2600
rect 450 2015 465 2585
rect 485 2015 500 2585
rect 450 2000 500 2015
rect 550 2585 600 2600
rect 550 2015 565 2585
rect 585 2015 600 2585
rect 550 2000 600 2015
rect 650 2585 700 2600
rect 650 2015 665 2585
rect 685 2015 700 2585
rect 650 2000 700 2015
rect 750 2585 800 2600
rect 750 2015 765 2585
rect 785 2015 800 2585
rect 750 2000 800 2015
rect 850 2585 900 2600
rect 850 2015 865 2585
rect 885 2015 900 2585
rect 850 2000 900 2015
rect 950 2585 1000 2600
rect 950 2015 965 2585
rect 985 2015 1000 2585
rect 950 2000 1000 2015
rect 1050 2585 1100 2600
rect 1050 2015 1065 2585
rect 1085 2015 1100 2585
rect 1050 2000 1100 2015
rect 1150 2585 1200 2600
rect 1250 2585 1300 2600
rect 1150 2015 1165 2585
rect 1185 2015 1200 2585
rect 1250 2015 1265 2585
rect 1285 2015 1300 2585
rect 1150 2000 1200 2015
rect 1250 2000 1300 2015
rect 1350 2585 1400 2600
rect 1350 2015 1365 2585
rect 1385 2015 1400 2585
rect 1350 2000 1400 2015
rect 1450 2585 1500 2600
rect 1450 2015 1465 2585
rect 1485 2015 1500 2585
rect 1450 2000 1500 2015
rect 1550 2585 1600 2600
rect 1550 2015 1565 2585
rect 1585 2015 1600 2585
rect 1550 2000 1600 2015
rect 1650 2585 1700 2600
rect 1650 2015 1665 2585
rect 1685 2015 1700 2585
rect 1650 2000 1700 2015
rect -145 1675 -95 1690
rect -145 1105 -130 1675
rect -110 1105 -95 1675
rect -145 1090 -95 1105
rect -45 1675 0 1690
rect -45 1105 -35 1675
rect -15 1105 0 1675
rect -45 1090 0 1105
rect 50 1675 100 1690
rect 50 1105 65 1675
rect 85 1105 100 1675
rect 50 1090 100 1105
rect 150 1675 200 1690
rect 150 1105 165 1675
rect 185 1105 200 1675
rect 150 1090 200 1105
rect 250 1675 300 1690
rect 350 1675 400 1690
rect 250 1105 265 1675
rect 285 1105 300 1675
rect 350 1105 365 1675
rect 385 1105 400 1675
rect 250 1090 300 1105
rect 350 1090 400 1105
rect 450 1675 500 1690
rect 450 1105 465 1675
rect 485 1105 500 1675
rect 450 1090 500 1105
rect 550 1675 600 1690
rect 550 1105 565 1675
rect 585 1105 600 1675
rect 550 1090 600 1105
rect 650 1675 700 1690
rect 650 1105 665 1675
rect 685 1105 700 1675
rect 650 1090 700 1105
rect 750 1675 800 1690
rect 750 1105 765 1675
rect 785 1105 800 1675
rect 750 1090 800 1105
rect 850 1675 900 1690
rect 850 1105 865 1675
rect 885 1105 900 1675
rect 850 1090 900 1105
rect 950 1675 1000 1690
rect 950 1105 965 1675
rect 985 1105 1000 1675
rect 950 1090 1000 1105
rect 1050 1675 1100 1690
rect 1050 1105 1065 1675
rect 1085 1105 1100 1675
rect 1050 1090 1100 1105
rect 1150 1675 1200 1690
rect 1250 1675 1300 1690
rect 1150 1105 1165 1675
rect 1185 1105 1200 1675
rect 1250 1105 1265 1675
rect 1285 1105 1300 1675
rect 1150 1090 1200 1105
rect 1250 1090 1300 1105
rect 1350 1675 1400 1690
rect 1350 1105 1365 1675
rect 1385 1105 1400 1675
rect 1350 1090 1400 1105
rect 1450 1675 1500 1690
rect 1450 1105 1465 1675
rect 1485 1105 1500 1675
rect 1450 1090 1500 1105
rect 1550 1675 1595 1690
rect 1550 1105 1565 1675
rect 1585 1105 1595 1675
rect 1550 1090 1595 1105
rect 1645 1675 1695 1690
rect 1645 1105 1660 1675
rect 1680 1105 1695 1675
rect 1645 1090 1695 1105
<< ndiffc >>
rect -135 280 -115 850
rect -35 280 -15 850
rect 65 280 85 850
rect 165 280 185 850
rect 265 280 285 850
rect 365 280 385 850
rect 465 280 485 850
rect 565 280 585 850
rect 665 280 685 850
rect 765 280 785 850
rect 865 280 885 850
rect 965 280 985 850
rect 1065 280 1085 850
rect 1165 280 1185 850
rect 1265 280 1285 850
rect 1365 280 1385 850
rect 1465 280 1485 850
rect 1565 280 1585 850
rect 1665 280 1685 850
<< pdiffc >>
rect -135 2015 -115 2585
rect -35 2015 -15 2585
rect 65 2015 85 2585
rect 165 2015 185 2585
rect 265 2015 285 2585
rect 365 2015 385 2585
rect 465 2015 485 2585
rect 565 2015 585 2585
rect 665 2015 685 2585
rect 765 2015 785 2585
rect 865 2015 885 2585
rect 965 2015 985 2585
rect 1065 2015 1085 2585
rect 1165 2015 1185 2585
rect 1265 2015 1285 2585
rect 1365 2015 1385 2585
rect 1465 2015 1485 2585
rect 1565 2015 1585 2585
rect 1665 2015 1685 2585
rect -130 1105 -110 1675
rect -35 1105 -15 1675
rect 65 1105 85 1675
rect 165 1105 185 1675
rect 265 1105 285 1675
rect 365 1105 385 1675
rect 465 1105 485 1675
rect 565 1105 585 1675
rect 665 1105 685 1675
rect 765 1105 785 1675
rect 865 1105 885 1675
rect 965 1105 985 1675
rect 1065 1105 1085 1675
rect 1165 1105 1185 1675
rect 1265 1105 1285 1675
rect 1365 1105 1385 1675
rect 1465 1105 1485 1675
rect 1565 1105 1585 1675
rect 1660 1105 1680 1675
<< psubdiff >>
rect 300 850 350 865
rect 300 280 315 850
rect 335 280 350 850
rect 300 265 350 280
rect 1200 850 1250 865
rect 1200 280 1215 850
rect 1235 280 1250 850
rect 1200 265 1250 280
<< nsubdiff >>
rect 300 2585 350 2600
rect 300 2015 315 2585
rect 335 2015 350 2585
rect 300 2000 350 2015
rect 1200 2585 1250 2600
rect 1200 2015 1215 2585
rect 1235 2015 1250 2585
rect 1200 2000 1250 2015
rect 300 1675 350 1690
rect 300 1105 315 1675
rect 335 1105 350 1675
rect 300 1090 350 1105
rect 1200 1675 1250 1690
rect 1200 1105 1215 1675
rect 1235 1105 1250 1675
rect 1200 1090 1250 1105
<< psubdiffcont >>
rect 315 280 335 850
rect 1215 280 1235 850
<< nsubdiffcont >>
rect 315 2015 335 2585
rect 1215 2015 1235 2585
rect 315 1105 335 1675
rect 1215 1105 1235 1675
<< poly >>
rect 0 2700 50 2715
rect 0 2680 15 2700
rect 35 2680 50 2700
rect -100 2645 -50 2660
rect -100 2625 -85 2645
rect -65 2625 -50 2645
rect -100 2600 -50 2625
rect 0 2600 50 2680
rect 600 2700 650 2715
rect 600 2680 615 2700
rect 635 2680 650 2700
rect 200 2645 250 2660
rect 200 2625 215 2645
rect 235 2625 250 2645
rect 100 2600 150 2620
rect 200 2600 250 2625
rect 400 2645 450 2660
rect 400 2625 415 2645
rect 435 2625 450 2645
rect 400 2600 450 2625
rect 500 2600 550 2620
rect 600 2600 650 2680
rect 900 2700 950 2715
rect 900 2680 915 2700
rect 935 2680 950 2700
rect 700 2645 750 2660
rect 700 2625 715 2645
rect 735 2625 750 2645
rect 700 2600 750 2625
rect 800 2645 850 2660
rect 800 2625 815 2645
rect 835 2625 850 2645
rect 800 2600 850 2625
rect 900 2600 950 2680
rect 1500 2700 1550 2715
rect 1500 2680 1515 2700
rect 1535 2680 1550 2700
rect 1100 2645 1150 2660
rect 1100 2625 1115 2645
rect 1135 2625 1150 2645
rect 1000 2600 1050 2620
rect 1100 2600 1150 2625
rect 1300 2645 1350 2660
rect 1300 2625 1315 2645
rect 1335 2625 1350 2645
rect 1300 2600 1350 2625
rect 1400 2600 1450 2620
rect 1500 2600 1550 2680
rect 1600 2645 1650 2660
rect 1600 2625 1615 2645
rect 1635 2625 1650 2645
rect 1600 2600 1650 2625
rect -100 1985 -50 2000
rect 0 1985 50 2000
rect 100 1965 150 2000
rect 200 1985 250 2000
rect 400 1985 450 2000
rect 100 1945 115 1965
rect 135 1945 150 1965
rect 100 1930 150 1945
rect 500 1965 550 2000
rect 600 1985 650 2000
rect 700 1985 750 2000
rect 800 1985 850 2000
rect 900 1985 950 2000
rect 500 1945 515 1965
rect 535 1945 550 1965
rect 500 1930 550 1945
rect 1000 1965 1050 2000
rect 1100 1985 1150 2000
rect 1300 1985 1350 2000
rect 1000 1945 1015 1965
rect 1035 1945 1050 1965
rect 1000 1930 1050 1945
rect 1400 1965 1450 2000
rect 1500 1985 1550 2000
rect 1600 1985 1650 2000
rect 1400 1945 1415 1965
rect 1435 1945 1450 1965
rect 1400 1930 1450 1945
rect 600 1855 650 1870
rect 600 1835 615 1855
rect 635 1835 650 1855
rect 0 1800 50 1815
rect 0 1780 15 1800
rect 35 1780 50 1800
rect -95 1735 -45 1750
rect -95 1715 -80 1735
rect -60 1715 -45 1735
rect -95 1690 -45 1715
rect 0 1690 50 1780
rect 100 1745 150 1760
rect 100 1725 115 1745
rect 135 1725 150 1745
rect 100 1690 150 1725
rect 200 1745 250 1760
rect 200 1725 215 1745
rect 235 1725 250 1745
rect 200 1690 250 1725
rect 400 1745 450 1760
rect 400 1725 415 1745
rect 435 1725 450 1745
rect 400 1690 450 1725
rect 500 1745 550 1760
rect 500 1725 515 1745
rect 535 1725 550 1745
rect 500 1690 550 1725
rect 600 1690 650 1835
rect 900 1855 950 1870
rect 900 1835 915 1855
rect 935 1835 950 1855
rect 700 1690 750 1705
rect 800 1690 850 1705
rect 900 1690 950 1835
rect 1500 1800 1550 1815
rect 1500 1780 1515 1800
rect 1535 1780 1550 1800
rect 1000 1745 1050 1760
rect 1000 1725 1015 1745
rect 1035 1725 1050 1745
rect 1000 1690 1050 1725
rect 1100 1745 1150 1760
rect 1100 1725 1115 1745
rect 1135 1725 1150 1745
rect 1100 1690 1150 1725
rect 1300 1745 1350 1760
rect 1300 1725 1315 1745
rect 1335 1725 1350 1745
rect 1300 1690 1350 1725
rect 1400 1745 1450 1760
rect 1400 1725 1415 1745
rect 1435 1725 1450 1745
rect 1400 1690 1450 1725
rect 1500 1690 1550 1780
rect 1595 1735 1645 1750
rect 1595 1715 1610 1735
rect 1630 1715 1645 1735
rect 1595 1690 1645 1715
rect -95 1075 -45 1090
rect 0 1075 50 1090
rect 100 1075 150 1090
rect 200 1075 250 1090
rect 400 1075 450 1090
rect 500 1075 550 1090
rect 600 1075 650 1090
rect 700 1075 750 1090
rect 800 1075 850 1090
rect 900 1075 950 1090
rect 1000 1075 1050 1090
rect 1100 1075 1150 1090
rect 1300 1075 1350 1090
rect 1400 1075 1450 1090
rect 1500 1075 1550 1090
rect 1595 1075 1645 1090
rect 700 1060 850 1075
rect 700 1040 765 1060
rect 785 1040 850 1060
rect 700 1025 850 1040
rect 200 905 250 920
rect 200 885 215 905
rect 235 885 250 905
rect -100 865 -50 880
rect 0 865 50 880
rect 100 865 150 880
rect 200 865 250 885
rect 400 905 450 920
rect 400 885 415 905
rect 435 885 450 905
rect 400 865 450 885
rect 1100 905 1150 920
rect 1100 885 1115 905
rect 1135 885 1150 905
rect 500 865 550 880
rect 600 865 650 880
rect 700 865 750 880
rect 800 865 850 880
rect 900 865 950 880
rect 1000 865 1050 880
rect 1100 865 1150 885
rect 1300 905 1350 920
rect 1300 885 1315 905
rect 1335 885 1350 905
rect 1300 865 1350 885
rect 1400 865 1450 880
rect 1500 865 1550 880
rect 1600 865 1650 880
rect -100 245 -50 265
rect -100 225 -85 245
rect -65 225 -50 245
rect -100 210 -50 225
rect 0 175 50 265
rect 100 230 150 265
rect 200 250 250 265
rect 400 250 450 265
rect 100 210 115 230
rect 135 210 150 230
rect 100 195 150 210
rect 500 230 550 265
rect 500 210 515 230
rect 535 210 550 230
rect 500 195 550 210
rect 0 155 15 175
rect 35 155 50 175
rect 0 140 50 155
rect 600 175 650 265
rect 700 245 750 265
rect 700 225 715 245
rect 735 225 750 245
rect 700 210 750 225
rect 800 245 850 265
rect 800 225 815 245
rect 835 225 850 245
rect 800 210 850 225
rect 600 155 615 175
rect 635 155 650 175
rect 600 140 650 155
rect 900 175 950 265
rect 1000 230 1050 265
rect 1100 250 1150 265
rect 1300 250 1350 265
rect 1000 210 1015 230
rect 1035 210 1050 230
rect 1000 195 1050 210
rect 1400 230 1450 265
rect 1400 210 1415 230
rect 1435 210 1450 230
rect 1400 195 1450 210
rect 900 155 915 175
rect 935 155 950 175
rect 900 140 950 155
rect 1500 175 1550 265
rect 1600 245 1650 265
rect 1600 225 1615 245
rect 1635 225 1650 245
rect 1600 210 1650 225
rect 1500 155 1515 175
rect 1535 155 1550 175
rect 1500 140 1550 155
<< polycont >>
rect 15 2680 35 2700
rect -85 2625 -65 2645
rect 615 2680 635 2700
rect 215 2625 235 2645
rect 415 2625 435 2645
rect 915 2680 935 2700
rect 715 2625 735 2645
rect 815 2625 835 2645
rect 1515 2680 1535 2700
rect 1115 2625 1135 2645
rect 1315 2625 1335 2645
rect 1615 2625 1635 2645
rect 115 1945 135 1965
rect 515 1945 535 1965
rect 1015 1945 1035 1965
rect 1415 1945 1435 1965
rect 615 1835 635 1855
rect 15 1780 35 1800
rect -80 1715 -60 1735
rect 115 1725 135 1745
rect 215 1725 235 1745
rect 415 1725 435 1745
rect 515 1725 535 1745
rect 915 1835 935 1855
rect 1515 1780 1535 1800
rect 1015 1725 1035 1745
rect 1115 1725 1135 1745
rect 1315 1725 1335 1745
rect 1415 1725 1435 1745
rect 1610 1715 1630 1735
rect 765 1040 785 1060
rect 215 885 235 905
rect 415 885 435 905
rect 1115 885 1135 905
rect 1315 885 1335 905
rect -85 225 -65 245
rect 115 210 135 230
rect 515 210 535 230
rect 15 155 35 175
rect 715 225 735 245
rect 815 225 835 245
rect 615 155 635 175
rect 1015 210 1035 230
rect 1415 210 1435 230
rect 915 155 935 175
rect 1615 225 1635 245
rect 1515 155 1535 175
<< locali >>
rect 5 2700 45 2710
rect 5 2680 15 2700
rect 35 2680 45 2700
rect 5 2670 45 2680
rect 605 2700 645 2710
rect 605 2680 615 2700
rect 635 2680 645 2700
rect 605 2670 645 2680
rect 905 2700 945 2710
rect 905 2680 915 2700
rect 935 2680 945 2700
rect 905 2670 945 2680
rect 1505 2700 1545 2710
rect 1505 2680 1515 2700
rect 1535 2680 1545 2700
rect 1505 2670 1545 2680
rect -145 2645 -55 2655
rect -145 2625 -85 2645
rect -65 2625 -55 2645
rect -145 2615 -55 2625
rect 155 2645 295 2655
rect 155 2625 215 2645
rect 235 2625 295 2645
rect 155 2615 295 2625
rect -145 2585 -105 2615
rect -145 2045 -135 2585
rect -150 2015 -135 2045
rect -115 2015 -105 2585
rect -150 2005 -105 2015
rect -45 2585 -5 2595
rect -45 2015 -35 2585
rect -15 2015 -5 2585
rect -205 1965 -165 1975
rect -205 1945 -195 1965
rect -175 1945 -165 1965
rect -205 940 -165 1945
rect -45 1965 -5 2015
rect 55 2585 95 2595
rect 55 2015 65 2585
rect 85 2015 95 2585
rect 55 2005 95 2015
rect 155 2585 195 2615
rect 155 2015 165 2585
rect 185 2015 195 2585
rect 155 2005 195 2015
rect 255 2595 295 2615
rect 355 2645 495 2655
rect 355 2625 415 2645
rect 435 2625 495 2645
rect 355 2615 495 2625
rect 355 2595 395 2615
rect 255 2585 395 2595
rect 255 2015 265 2585
rect 285 2015 315 2585
rect 335 2015 365 2585
rect 385 2015 395 2585
rect 255 2005 395 2015
rect 455 2585 495 2615
rect 655 2645 895 2655
rect 655 2625 715 2645
rect 735 2625 815 2645
rect 835 2625 895 2645
rect 655 2615 895 2625
rect 455 2015 465 2585
rect 485 2015 495 2585
rect 455 2005 495 2015
rect 555 2585 595 2595
rect 555 2015 565 2585
rect 585 2015 595 2585
rect 555 2005 595 2015
rect 655 2585 695 2615
rect 655 2015 665 2585
rect 685 2015 695 2585
rect -45 1945 -35 1965
rect -15 1945 -5 1965
rect -45 1935 -5 1945
rect 105 1965 145 1975
rect 105 1945 115 1965
rect 135 1945 145 1965
rect 105 1935 145 1945
rect 5 1800 45 1810
rect 5 1780 15 1800
rect 35 1780 45 1800
rect 5 1770 45 1780
rect 105 1745 145 1755
rect -140 1735 -50 1745
rect -140 1715 -80 1735
rect -60 1715 -50 1735
rect 105 1725 115 1745
rect 135 1725 145 1745
rect 105 1715 145 1725
rect 205 1745 245 1755
rect 205 1725 215 1745
rect 235 1725 245 1745
rect 205 1715 245 1725
rect -140 1705 -50 1715
rect -140 1675 -100 1705
rect 265 1685 385 2005
rect 505 1965 545 1975
rect 505 1945 515 1965
rect 535 1945 545 1965
rect 505 1935 545 1945
rect 655 1920 695 2015
rect 755 2585 795 2615
rect 755 2015 765 2585
rect 785 2015 795 2585
rect 755 1985 795 2015
rect 855 2585 895 2615
rect 1055 2645 1195 2655
rect 1055 2625 1115 2645
rect 1135 2625 1195 2645
rect 1055 2615 1195 2625
rect 855 2015 865 2585
rect 885 2015 895 2585
rect 855 1920 895 2015
rect 955 2585 995 2595
rect 955 2015 965 2585
rect 985 2015 995 2585
rect 955 2005 995 2015
rect 1055 2585 1095 2615
rect 1055 2015 1065 2585
rect 1085 2015 1095 2585
rect 1055 2005 1095 2015
rect 1155 2595 1195 2615
rect 1255 2645 1395 2655
rect 1255 2625 1315 2645
rect 1335 2625 1395 2645
rect 1255 2615 1395 2625
rect 1605 2645 1695 2655
rect 1605 2625 1615 2645
rect 1635 2625 1695 2645
rect 1605 2615 1695 2625
rect 1255 2595 1295 2615
rect 1155 2585 1295 2595
rect 1155 2015 1165 2585
rect 1185 2015 1215 2585
rect 1235 2015 1265 2585
rect 1285 2015 1295 2585
rect 1155 2005 1295 2015
rect 1355 2585 1395 2615
rect 1355 2015 1365 2585
rect 1385 2015 1395 2585
rect 1355 2005 1395 2015
rect 1455 2585 1495 2595
rect 1455 2015 1465 2585
rect 1485 2015 1495 2585
rect 1455 2005 1495 2015
rect 1555 2585 1595 2595
rect 1555 2015 1565 2585
rect 1585 2015 1595 2585
rect 1005 1965 1045 1975
rect 1005 1945 1015 1965
rect 1035 1945 1045 1965
rect 1005 1935 1045 1945
rect 655 1910 735 1920
rect 655 1890 665 1910
rect 685 1890 735 1910
rect 655 1880 735 1890
rect 605 1855 645 1865
rect 605 1835 615 1855
rect 635 1835 645 1855
rect 605 1825 645 1835
rect 405 1745 445 1755
rect 405 1725 415 1745
rect 435 1725 445 1745
rect 405 1715 445 1725
rect 505 1745 545 1755
rect 505 1725 515 1745
rect 535 1725 545 1745
rect 505 1715 545 1725
rect -140 1135 -130 1675
rect -145 1105 -130 1135
rect -110 1105 -100 1675
rect -145 1095 -100 1105
rect -45 1675 -5 1685
rect -45 1105 -35 1675
rect -15 1105 -5 1675
rect -45 1000 -5 1105
rect 55 1675 95 1685
rect 55 1105 65 1675
rect 85 1105 95 1675
rect 55 1075 95 1105
rect 155 1675 195 1685
rect 155 1105 165 1675
rect 185 1105 195 1675
rect 155 1095 195 1105
rect 255 1675 395 1685
rect 255 1105 265 1675
rect 285 1105 315 1675
rect 335 1105 365 1675
rect 385 1105 395 1675
rect 255 1095 395 1105
rect 455 1675 495 1685
rect 455 1105 465 1675
rect 485 1105 495 1675
rect 455 1095 495 1105
rect 555 1675 595 1685
rect 555 1105 565 1675
rect 585 1105 595 1675
rect 555 1075 595 1105
rect 55 1035 595 1075
rect 655 1675 695 1685
rect 655 1105 665 1675
rect 685 1105 695 1675
rect 655 1015 695 1105
rect -45 960 95 1000
rect -205 900 -5 940
rect -145 850 -105 860
rect -145 280 -135 850
rect -115 280 -105 850
rect -145 255 -105 280
rect -45 850 -5 900
rect -45 280 -35 850
rect -15 280 -5 850
rect -45 270 -5 280
rect 55 850 95 960
rect 555 975 695 1015
rect 55 280 65 850
rect 85 280 95 850
rect 55 270 95 280
rect 155 905 295 915
rect 155 885 215 905
rect 235 885 295 905
rect 155 875 295 885
rect 155 850 195 875
rect 155 280 165 850
rect 185 280 195 850
rect 155 270 195 280
rect 255 865 295 875
rect 355 905 495 915
rect 355 885 415 905
rect 435 885 495 905
rect 355 875 495 885
rect 255 860 300 865
rect 355 860 395 875
rect 255 850 395 860
rect 255 280 265 850
rect 285 280 315 850
rect 335 280 365 850
rect 385 280 395 850
rect 255 270 395 280
rect 455 850 495 875
rect 455 280 465 850
rect 485 280 495 850
rect 455 270 495 280
rect 555 850 595 975
rect 715 955 735 1880
rect 815 1910 895 1920
rect 815 1890 865 1910
rect 885 1890 895 1910
rect 815 1880 895 1890
rect 755 1675 795 1705
rect 755 1105 765 1675
rect 785 1105 795 1675
rect 755 1060 795 1105
rect 755 1040 765 1060
rect 785 1040 795 1060
rect 755 1030 795 1040
rect 555 280 565 850
rect 585 280 595 850
rect 555 270 595 280
rect 655 915 735 955
rect 815 955 835 1880
rect 905 1855 945 1865
rect 905 1835 915 1855
rect 935 1835 945 1855
rect 905 1825 945 1835
rect 1005 1745 1045 1755
rect 1005 1725 1015 1745
rect 1035 1725 1045 1745
rect 1005 1715 1045 1725
rect 1105 1745 1145 1755
rect 1105 1725 1115 1745
rect 1135 1725 1145 1745
rect 1105 1715 1145 1725
rect 1165 1685 1285 2005
rect 1405 1965 1445 1975
rect 1405 1945 1415 1965
rect 1435 1945 1445 1965
rect 1405 1935 1445 1945
rect 1555 1965 1595 2015
rect 1655 2585 1695 2615
rect 1655 2015 1665 2585
rect 1685 2045 1695 2585
rect 1685 2015 1700 2045
rect 1655 2005 1700 2015
rect 1555 1945 1565 1965
rect 1585 1945 1595 1965
rect 1555 1935 1595 1945
rect 1715 1965 1755 1975
rect 1715 1945 1725 1965
rect 1745 1945 1755 1965
rect 1505 1800 1545 1810
rect 1505 1780 1515 1800
rect 1535 1780 1545 1800
rect 1505 1770 1545 1780
rect 1305 1745 1345 1755
rect 1305 1725 1315 1745
rect 1335 1725 1345 1745
rect 1305 1715 1345 1725
rect 1405 1745 1445 1755
rect 1405 1725 1415 1745
rect 1435 1725 1445 1745
rect 1405 1715 1445 1725
rect 1600 1735 1690 1745
rect 1600 1715 1610 1735
rect 1630 1715 1690 1735
rect 1600 1705 1690 1715
rect 855 1675 895 1685
rect 855 1105 865 1675
rect 885 1105 895 1675
rect 855 1015 895 1105
rect 955 1675 995 1685
rect 955 1105 965 1675
rect 985 1105 995 1675
rect 955 1075 995 1105
rect 1055 1675 1095 1685
rect 1055 1105 1065 1675
rect 1085 1105 1095 1675
rect 1055 1095 1095 1105
rect 1155 1675 1295 1685
rect 1155 1105 1165 1675
rect 1185 1105 1215 1675
rect 1235 1105 1265 1675
rect 1285 1105 1295 1675
rect 1155 1095 1295 1105
rect 1355 1675 1395 1685
rect 1355 1105 1365 1675
rect 1385 1105 1395 1675
rect 1355 1095 1395 1105
rect 1455 1675 1495 1685
rect 1455 1105 1465 1675
rect 1485 1105 1495 1675
rect 1455 1075 1495 1105
rect 955 1035 1495 1075
rect 1555 1675 1595 1685
rect 1555 1105 1565 1675
rect 1585 1105 1595 1675
rect 855 975 995 1015
rect 1555 1000 1595 1105
rect 1650 1675 1690 1705
rect 1650 1105 1660 1675
rect 1680 1135 1690 1675
rect 1680 1105 1695 1135
rect 1650 1095 1695 1105
rect 815 915 895 955
rect 655 850 695 915
rect 655 280 665 850
rect 685 280 695 850
rect 655 255 695 280
rect 755 850 795 860
rect 755 280 765 850
rect 785 280 795 850
rect 755 255 795 280
rect 855 850 895 915
rect 855 280 865 850
rect 885 280 895 850
rect 855 255 895 280
rect 955 850 995 975
rect 1455 960 1595 1000
rect 955 280 965 850
rect 985 280 995 850
rect 955 270 995 280
rect 1055 905 1195 915
rect 1055 885 1115 905
rect 1135 885 1195 905
rect 1055 875 1195 885
rect 1055 850 1095 875
rect 1055 280 1065 850
rect 1085 280 1095 850
rect 1055 270 1095 280
rect 1155 860 1195 875
rect 1255 905 1395 915
rect 1255 885 1315 905
rect 1335 885 1395 905
rect 1255 875 1395 885
rect 1255 865 1295 875
rect 1250 860 1295 865
rect 1155 850 1295 860
rect 1155 280 1165 850
rect 1185 280 1215 850
rect 1235 280 1265 850
rect 1285 280 1295 850
rect 1155 270 1295 280
rect 1355 850 1395 875
rect 1355 280 1365 850
rect 1385 280 1395 850
rect 1355 270 1395 280
rect 1455 850 1495 960
rect 1715 940 1755 1945
rect 1455 280 1465 850
rect 1485 280 1495 850
rect 1455 270 1495 280
rect 1555 900 1755 940
rect 1555 850 1595 900
rect 1555 280 1565 850
rect 1585 280 1595 850
rect 1555 270 1595 280
rect 1655 850 1695 860
rect 1655 280 1665 850
rect 1685 280 1695 850
rect 1655 255 1695 280
rect -145 245 -55 255
rect -145 225 -85 245
rect -65 225 -55 245
rect 655 245 895 255
rect -145 215 -55 225
rect 105 230 145 240
rect 105 210 115 230
rect 135 210 145 230
rect 105 200 145 210
rect 505 230 545 240
rect 505 210 515 230
rect 535 210 545 230
rect 655 225 715 245
rect 735 225 815 245
rect 835 225 895 245
rect 1605 245 1695 255
rect 655 215 895 225
rect 1005 230 1045 240
rect 505 200 545 210
rect 1005 210 1015 230
rect 1035 210 1045 230
rect 1005 200 1045 210
rect 1405 230 1445 240
rect 1405 210 1415 230
rect 1435 210 1445 230
rect 1605 225 1615 245
rect 1635 225 1695 245
rect 1605 215 1695 225
rect 1405 200 1445 210
rect 5 175 45 185
rect 5 155 15 175
rect 35 155 45 175
rect 5 145 45 155
rect 605 175 645 185
rect 605 155 615 175
rect 635 155 645 175
rect 605 145 645 155
rect 905 175 945 185
rect 905 155 915 175
rect 935 155 945 175
rect 905 145 945 155
rect 1505 175 1545 185
rect 1505 155 1515 175
rect 1535 155 1545 175
rect 1505 145 1545 155
<< viali >>
rect 15 2680 35 2700
rect 615 2680 635 2700
rect 915 2680 935 2700
rect 1515 2680 1535 2700
rect -135 2015 -115 2585
rect -195 1945 -175 1965
rect 165 2015 185 2585
rect 265 2015 285 2585
rect 315 2015 335 2585
rect 365 2015 385 2585
rect 465 2015 485 2585
rect -35 1945 -15 1965
rect 115 1945 135 1965
rect 15 1780 35 1800
rect 115 1725 135 1745
rect 215 1725 235 1745
rect 515 1945 535 1965
rect 1065 2015 1085 2585
rect 1165 2015 1185 2585
rect 1215 2015 1235 2585
rect 1265 2015 1285 2585
rect 1365 2015 1385 2585
rect 1015 1945 1035 1965
rect 665 1890 685 1910
rect 615 1835 635 1855
rect 415 1725 435 1745
rect 515 1725 535 1745
rect -130 1105 -110 1675
rect 265 1105 285 1675
rect 315 1105 335 1675
rect 365 1105 385 1675
rect -135 280 -115 850
rect 165 280 185 850
rect 265 280 285 850
rect 315 280 335 850
rect 365 280 385 850
rect 465 280 485 850
rect 865 1890 885 1910
rect 765 1105 785 1675
rect 915 1835 935 1855
rect 1015 1725 1035 1745
rect 1115 1725 1135 1745
rect 1415 1945 1435 1965
rect 1665 2015 1685 2585
rect 1565 1945 1585 1965
rect 1725 1945 1745 1965
rect 1515 1780 1535 1800
rect 1315 1725 1335 1745
rect 1415 1725 1435 1745
rect 1165 1105 1185 1675
rect 1215 1105 1235 1675
rect 1265 1105 1285 1675
rect 1660 1105 1680 1675
rect 1065 280 1085 850
rect 1165 280 1185 850
rect 1215 280 1235 850
rect 1265 280 1285 850
rect 1365 280 1385 850
rect 1665 280 1685 850
rect 115 210 135 230
rect 515 210 535 230
rect 1015 210 1035 230
rect 1415 210 1435 230
rect 15 155 35 175
rect 615 155 635 175
rect 915 155 935 175
rect 1515 155 1535 175
<< metal1 >>
rect -245 2700 1795 2710
rect -245 2680 15 2700
rect 35 2680 615 2700
rect 635 2680 915 2700
rect 935 2680 1515 2700
rect 1535 2680 1795 2700
rect -245 2670 1795 2680
rect -245 2585 1700 2595
rect -245 2015 -135 2585
rect -115 2015 165 2585
rect 185 2015 265 2585
rect 285 2015 315 2585
rect 335 2015 365 2585
rect 385 2015 465 2585
rect 485 2015 1065 2585
rect 1085 2015 1165 2585
rect 1185 2015 1215 2585
rect 1235 2015 1265 2585
rect 1285 2015 1365 2585
rect 1385 2015 1665 2585
rect 1685 2015 1700 2585
rect -245 2005 1700 2015
rect -205 1965 545 1975
rect -205 1945 -195 1965
rect -175 1945 -35 1965
rect -15 1945 115 1965
rect 135 1945 515 1965
rect 535 1945 545 1965
rect -205 1935 545 1945
rect 1005 1965 1755 1975
rect 1005 1945 1015 1965
rect 1035 1945 1415 1965
rect 1435 1945 1565 1965
rect 1585 1945 1725 1965
rect 1745 1945 1755 1965
rect 1005 1935 1755 1945
rect -245 1910 1755 1920
rect -245 1890 665 1910
rect 685 1890 865 1910
rect 885 1890 1755 1910
rect -245 1880 1755 1890
rect -245 1855 1755 1865
rect -245 1835 615 1855
rect 635 1835 915 1855
rect 935 1835 1755 1855
rect -245 1825 1755 1835
rect -245 1800 1755 1810
rect -245 1780 15 1800
rect 35 1780 1515 1800
rect 1535 1780 1755 1800
rect -245 1770 1755 1780
rect -245 1745 1755 1755
rect -245 1725 115 1745
rect 135 1725 215 1745
rect 235 1725 415 1745
rect 435 1725 515 1745
rect 535 1725 1015 1745
rect 1035 1725 1115 1745
rect 1135 1725 1315 1745
rect 1335 1725 1415 1745
rect 1435 1725 1755 1745
rect -245 1715 1755 1725
rect -245 1675 1695 1685
rect -245 1105 -130 1675
rect -110 1105 265 1675
rect 285 1105 315 1675
rect 335 1105 365 1675
rect 385 1105 765 1675
rect 785 1105 1165 1675
rect 1185 1105 1215 1675
rect 1235 1105 1265 1675
rect 1285 1105 1660 1675
rect 1680 1105 1695 1675
rect -245 1095 1695 1105
rect -245 850 1700 860
rect -245 280 -135 850
rect -115 280 165 850
rect 185 280 265 850
rect 285 280 315 850
rect 335 280 365 850
rect 385 280 465 850
rect 485 280 1065 850
rect 1085 280 1165 850
rect 1185 280 1215 850
rect 1235 280 1265 850
rect 1285 280 1365 850
rect 1385 280 1665 850
rect 1685 280 1700 850
rect -245 270 1700 280
rect -245 230 1695 240
rect -245 210 115 230
rect 135 210 515 230
rect 535 210 1015 230
rect 1035 210 1415 230
rect 1435 210 1695 230
rect -245 200 1695 210
rect -245 175 1690 185
rect -245 155 15 175
rect 35 155 615 175
rect 635 155 915 175
rect 935 155 1515 175
rect 1535 155 1690 175
rect -245 145 1690 155
<< labels >>
rlabel metal1 -245 2670 -205 2710 7 vcp
rlabel metal1 -245 2005 -205 2595 7 VDD
rlabel metal1 -245 270 -205 860 7 GND
rlabel metal1 -245 1095 -205 1685 7 VDD
rlabel metal1 -245 200 -205 240 7 vbn
rlabel metal1 -245 145 -205 185 7 vcn
rlabel metal1 -245 1880 -205 1920 7 vout
rlabel metal1 -245 1825 -205 1865 7 v2
rlabel metal1 -245 1770 -205 1810 7 v1
rlabel metal1 -245 1715 -205 1755 7 vbp
rlabel locali 65 1105 85 1675 1 net4
rlabel locali 165 1105 185 1675 1 net7
rlabel locali 465 1105 485 1675 1 net8
rlabel locali 665 1105 685 1675 1 net6
rlabel locali 565 2015 585 2585 1 net3
rlabel locali 65 2015 85 2585 1 net2
rlabel locali -35 2015 -15 2585 1 net1
rlabel locali -35 1105 -15 1675 1 net5
rlabel locali 1465 280 1485 850 1 net11
rlabel locali 1065 1105 1085 1675 1 net14
<< end >>
