magic
tech sky130A
timestamp 1614270932
use inverter_ports  inverter_ports_0
timestamp 1614270859
transform 1 0 35 0 1 365
box -215 -55 -50 860
use dff_4_wide_ports  dff_4_wide_ports_3
timestamp 1614264236
transform 1 0 730 0 1 -105
box -60 95 265 1330
use dff_4_wide_ports  dff_4_wide_ports_2
timestamp 1614264236
transform 1 0 495 0 1 -105
box -60 95 265 1330
use dff_4_wide_ports  dff_4_wide_ports_1
timestamp 1614264236
transform 1 0 260 0 1 -105
box -60 95 265 1330
use dff_4_wide_ports  dff_4_wide_ports_0
timestamp 1614264236
transform 1 0 25 0 1 -105
box -60 95 265 1330
<< end >>
