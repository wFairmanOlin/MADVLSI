magic
tech sky130A
timestamp 1614184383
<< nwell >>
rect -155 730 265 1280
<< nmos >>
rect 10 595 25 695
rect 50 595 65 695
rect 115 595 130 695
rect 180 595 195 695
rect 10 225 25 325
rect 50 225 65 325
rect 115 225 130 325
rect 180 225 195 325
<< pmos >>
rect 10 1115 25 1215
rect 75 1115 90 1215
rect 140 1115 155 1215
rect 180 1115 195 1215
rect 10 765 25 865
rect 75 765 90 865
rect 140 765 155 865
rect 180 765 195 865
<< ndiff >>
rect -40 680 10 695
rect -40 610 -25 680
rect -5 610 10 680
rect -40 595 10 610
rect 25 595 50 695
rect 65 680 115 695
rect 65 610 80 680
rect 100 610 115 680
rect 65 595 115 610
rect 130 680 180 695
rect 130 610 145 680
rect 165 610 180 680
rect 130 595 180 610
rect 195 680 245 695
rect 195 610 210 680
rect 230 610 245 680
rect 195 595 245 610
rect -40 310 10 325
rect -40 240 -25 310
rect -5 240 10 310
rect -40 225 10 240
rect 25 225 50 325
rect 65 310 115 325
rect 65 240 80 310
rect 100 240 115 310
rect 65 225 115 240
rect 130 310 180 325
rect 130 240 145 310
rect 165 240 180 310
rect 130 225 180 240
rect 195 310 245 325
rect 195 240 210 310
rect 230 240 245 310
rect 195 225 245 240
<< pdiff >>
rect -40 1200 10 1215
rect -40 1130 -25 1200
rect -5 1130 10 1200
rect -40 1115 10 1130
rect 25 1200 75 1215
rect 25 1130 40 1200
rect 60 1130 75 1200
rect 25 1115 75 1130
rect 90 1200 140 1215
rect 90 1130 105 1200
rect 125 1130 140 1200
rect 90 1115 140 1130
rect 155 1115 180 1215
rect 195 1200 245 1215
rect 195 1130 210 1200
rect 230 1130 245 1200
rect 195 1115 245 1130
rect -40 850 10 865
rect -40 780 -25 850
rect -5 780 10 850
rect -40 765 10 780
rect 25 850 75 865
rect 25 780 40 850
rect 60 780 75 850
rect 25 765 75 780
rect 90 850 140 865
rect 90 780 105 850
rect 125 780 140 850
rect 90 765 140 780
rect 155 765 180 865
rect 195 850 245 865
rect 195 780 210 850
rect 230 780 245 850
rect 195 765 245 780
<< ndiffc >>
rect -25 610 -5 680
rect 80 610 100 680
rect 145 610 165 680
rect 210 610 230 680
rect -25 240 -5 310
rect 80 240 100 310
rect 145 240 165 310
rect 210 240 230 310
<< pdiffc >>
rect -25 1130 -5 1200
rect 40 1130 60 1200
rect 105 1130 125 1200
rect 210 1130 230 1200
rect -25 780 -5 850
rect 40 780 60 850
rect 105 780 125 850
rect 210 780 230 850
<< psubdiff >>
rect -145 490 -95 505
rect -145 420 -130 490
rect -110 420 -95 490
rect -145 405 -95 420
<< nsubdiff >>
rect -120 850 -70 865
rect -120 780 -105 850
rect -85 780 -70 850
rect -120 765 -70 780
<< psubdiffcont >>
rect -130 420 -110 490
<< nsubdiffcont >>
rect -105 780 -85 850
<< poly >>
rect 10 1215 25 1230
rect 75 1215 90 1230
rect 140 1215 155 1230
rect 180 1215 195 1230
rect 10 1050 25 1115
rect 75 1060 90 1115
rect 75 1050 115 1060
rect 10 1035 35 1050
rect 20 950 35 1035
rect 75 1030 85 1050
rect 105 1030 115 1050
rect 75 1020 115 1030
rect 140 995 155 1115
rect 180 1020 195 1115
rect 180 1010 230 1020
rect 180 1005 200 1010
rect 10 935 35 950
rect 120 980 155 995
rect 190 990 200 1005
rect 220 990 230 1010
rect 190 980 230 990
rect 10 865 25 935
rect 50 910 90 920
rect 50 890 60 910
rect 80 890 90 910
rect 50 880 90 890
rect 75 865 90 880
rect 120 890 135 980
rect 160 945 200 955
rect 160 925 170 945
rect 190 925 200 945
rect 160 915 200 925
rect 120 875 155 890
rect 140 865 155 875
rect 180 865 195 915
rect 10 695 25 765
rect 75 750 90 765
rect 140 750 155 765
rect 50 735 90 750
rect 115 735 155 750
rect 50 695 65 735
rect 115 695 130 735
rect 180 695 195 765
rect 10 585 25 595
rect -5 570 25 585
rect -5 415 10 570
rect 50 540 65 595
rect 50 530 90 540
rect 50 510 60 530
rect 80 510 90 530
rect 50 500 90 510
rect 115 480 130 595
rect 35 465 75 475
rect 35 445 45 465
rect 65 445 75 465
rect 35 435 75 445
rect 100 465 130 480
rect -5 400 25 415
rect 10 325 25 400
rect 50 325 65 435
rect 100 385 115 465
rect 180 460 195 595
rect 165 445 195 460
rect 140 435 180 445
rect 140 415 150 435
rect 170 415 180 435
rect 140 405 180 415
rect 100 370 130 385
rect 115 325 130 370
rect 180 370 220 380
rect 180 350 190 370
rect 210 350 220 370
rect 180 340 220 350
rect 180 325 195 340
rect 10 210 25 225
rect 50 210 65 225
rect 115 210 130 225
rect 180 210 195 225
rect -15 200 25 210
rect -15 180 -5 200
rect 15 180 25 200
rect -15 170 25 180
rect 115 200 155 210
rect 115 180 125 200
rect 145 180 155 200
rect 115 170 155 180
<< polycont >>
rect 85 1030 105 1050
rect 200 990 220 1010
rect 60 890 80 910
rect 170 925 190 945
rect 60 510 80 530
rect 45 445 65 465
rect 150 415 170 435
rect 190 350 210 370
rect -5 180 15 200
rect 125 180 145 200
<< locali >>
rect -35 1200 5 1210
rect -35 1130 -25 1200
rect -5 1130 5 1200
rect -35 1120 5 1130
rect 30 1200 70 1210
rect 30 1130 40 1200
rect 60 1130 70 1200
rect 30 1120 70 1130
rect 95 1200 135 1210
rect 95 1130 105 1200
rect 125 1130 135 1200
rect 95 1120 135 1130
rect 200 1200 240 1210
rect 200 1130 210 1200
rect 230 1130 240 1200
rect 200 1120 240 1130
rect 35 920 55 1120
rect 200 1060 220 1120
rect 75 1050 115 1060
rect 75 1030 85 1050
rect 105 1040 115 1050
rect 150 1040 220 1060
rect 105 1030 130 1040
rect 75 1020 130 1030
rect 35 910 90 920
rect 35 900 60 910
rect 50 890 60 900
rect 80 890 90 910
rect 50 880 90 890
rect 110 860 130 1020
rect 150 955 170 1040
rect 190 1010 230 1020
rect 190 990 200 1010
rect 220 1000 230 1010
rect 220 990 240 1000
rect 190 980 240 990
rect 150 945 200 955
rect 150 925 170 945
rect 190 925 200 945
rect 150 915 200 925
rect 220 860 240 980
rect -115 850 -75 860
rect -115 780 -105 850
rect -85 780 -75 850
rect -115 770 -75 780
rect -35 850 5 860
rect -35 780 -25 850
rect -5 780 5 850
rect -35 770 5 780
rect 30 850 70 860
rect 30 780 40 850
rect 60 780 70 850
rect 30 770 70 780
rect 95 850 135 860
rect 95 780 105 850
rect 125 780 135 850
rect 95 770 135 780
rect 200 850 240 860
rect 200 780 210 850
rect 230 780 240 850
rect 200 770 240 780
rect 50 750 70 770
rect 200 750 220 770
rect 50 730 90 750
rect 70 690 90 730
rect 155 730 220 750
rect 155 690 175 730
rect -40 680 5 690
rect -40 610 -25 680
rect -5 610 5 680
rect -40 600 5 610
rect 70 680 110 690
rect 70 610 80 680
rect 100 610 110 680
rect 70 600 110 610
rect 135 680 175 690
rect 135 610 145 680
rect 165 610 175 680
rect 135 600 175 610
rect 200 680 240 690
rect 200 610 210 680
rect 230 610 240 680
rect 200 600 240 610
rect 70 580 90 600
rect 10 560 90 580
rect -140 490 -100 500
rect -140 420 -130 490
rect -110 420 -100 490
rect 10 475 30 560
rect 50 530 90 540
rect 50 510 60 530
rect 80 520 90 530
rect 80 510 115 520
rect 50 500 115 510
rect 10 465 75 475
rect 10 455 45 465
rect 35 445 45 455
rect 65 445 75 465
rect 35 435 75 445
rect -140 410 -100 420
rect 95 365 115 500
rect 155 485 175 600
rect 155 465 220 485
rect 90 345 115 365
rect 140 435 180 445
rect 140 415 150 435
rect 170 415 180 435
rect 140 405 180 415
rect 90 320 110 345
rect 140 320 160 405
rect 200 380 220 465
rect 180 370 220 380
rect 180 350 190 370
rect 210 350 220 370
rect 180 340 220 350
rect -40 310 5 320
rect -40 240 -25 310
rect -5 240 5 310
rect -40 230 5 240
rect 70 310 110 320
rect 70 240 80 310
rect 100 240 110 310
rect 70 230 110 240
rect 135 310 175 320
rect 135 240 145 310
rect 165 240 175 310
rect 135 230 175 240
rect 200 310 245 320
rect 200 240 210 310
rect 230 240 245 310
rect 200 230 245 240
rect -15 200 25 210
rect -15 190 -5 200
rect -40 180 -5 190
rect 15 190 25 200
rect 115 200 155 210
rect 115 190 125 200
rect 15 180 125 190
rect 145 190 155 200
rect 145 180 245 190
rect -40 170 245 180
<< end >>
