magic
tech sky130A
magscale 1 2
timestamp 1614019722
<< error_p >>
rect 85 1320 100 1720
rect 130 1320 154 1720
rect 215 1320 230 1365
<< nmos >>
rect 100 1120 130 1320
rect 230 1120 260 1320
rect 100 560 130 760
rect 230 560 260 760
rect 100 0 130 200
rect 230 0 260 200
<< ndiff >>
rect 0 1290 100 1720
rect 0 1150 30 1290
rect 70 1150 100 1290
rect 0 1120 100 1150
rect 130 1290 230 1720
rect 130 1150 160 1290
rect 200 1150 230 1290
rect 130 1120 230 1150
rect 260 1290 360 1320
rect 260 1150 290 1290
rect 330 1150 360 1290
rect 260 1120 360 1150
rect 0 730 100 760
rect 0 590 30 730
rect 70 590 100 730
rect 0 560 100 590
rect 130 730 230 760
rect 130 590 160 730
rect 200 590 230 730
rect 130 560 230 590
rect 260 730 360 760
rect 260 590 290 730
rect 330 590 360 730
rect 260 560 360 590
rect 0 170 100 200
rect 0 30 30 170
rect 70 30 100 170
rect 0 0 100 30
rect 130 170 230 200
rect 130 30 160 170
rect 200 30 230 170
rect 130 0 230 30
rect 260 170 360 200
rect 260 30 290 170
rect 330 30 360 170
rect 260 0 360 30
<< ndiffc >>
rect 30 1150 70 1290
rect 160 1150 200 1290
rect 290 1150 330 1290
rect 30 590 70 730
rect 160 590 200 730
rect 290 590 330 730
rect 30 30 70 170
rect 160 30 200 170
rect 290 30 330 170
<< psubdiff >>
rect -100 170 0 200
rect -100 30 -70 170
rect -20 30 0 170
rect -100 0 0 30
<< psubdiffcont >>
rect -70 30 -20 170
<< poly >>
rect 100 1320 130 1750
rect 230 1320 260 1350
rect 100 760 130 1120
rect 230 1090 260 1120
rect 230 760 260 790
rect 100 540 130 560
rect 0 510 130 540
rect 230 530 260 560
rect 230 510 310 530
rect 0 250 30 510
rect 230 470 250 510
rect 290 470 310 510
rect 100 440 180 460
rect 230 450 310 470
rect 100 400 120 440
rect 160 400 180 440
rect 100 380 180 400
rect 150 320 180 380
rect 150 290 260 320
rect 0 220 130 250
rect 100 200 130 220
rect 230 200 260 290
rect 100 -30 130 0
rect 230 -30 260 0
<< polycont >>
rect 250 470 290 510
rect 120 400 160 440
<< locali >>
rect 10 1290 90 1310
rect 10 1150 30 1290
rect 70 1150 90 1290
rect 10 1130 90 1150
rect 140 1290 220 1310
rect 140 1150 160 1290
rect 200 1150 220 1290
rect 140 1130 220 1150
rect 270 1290 350 1310
rect 270 1150 290 1290
rect 330 1150 350 1290
rect 270 1130 350 1150
rect 10 730 90 750
rect 10 590 30 730
rect 70 590 90 730
rect 10 570 90 590
rect 140 730 220 750
rect 140 590 160 730
rect 200 590 220 730
rect 140 570 220 590
rect 270 730 350 750
rect 270 590 290 730
rect 330 590 350 730
rect 270 570 350 590
rect 140 460 180 570
rect 100 440 180 460
rect 230 510 310 530
rect 230 470 250 510
rect 290 470 310 510
rect 230 450 310 470
rect 100 400 120 440
rect 160 400 180 440
rect 100 380 180 400
rect 270 270 310 450
rect 160 230 310 270
rect 160 190 200 230
rect -90 170 90 190
rect -90 30 -70 170
rect -20 30 30 170
rect 70 30 90 170
rect -90 10 90 30
rect 140 170 220 190
rect 140 30 160 170
rect 200 30 220 170
rect 140 10 220 30
rect 270 170 350 190
rect 270 30 290 170
rect 330 30 350 170
rect 270 10 350 30
<< end >>
