magic
tech sky130A
timestamp 1616129296
<< nwell >>
rect -95 1935 780 2695
rect -85 1660 770 1935
rect -85 955 760 1660
<< nmos >>
rect 0 0 50 600
rect 100 0 150 600
rect 200 0 250 600
rect 400 0 450 600
rect 500 0 550 600
rect 600 0 650 600
<< pmos >>
rect 0 2000 50 2600
rect 100 2000 150 2600
rect 200 2000 250 2600
rect 400 2000 450 2600
rect 500 2000 550 2600
rect 600 2000 650 2600
rect 0 1000 50 1600
rect 100 1000 150 1600
rect 200 1000 250 1600
rect 400 1000 450 1600
rect 500 1000 550 1600
rect 600 1000 650 1600
<< ndiff >>
rect -50 585 0 600
rect -50 15 -35 585
rect -15 15 0 585
rect -50 0 0 15
rect 50 585 100 600
rect 50 15 65 585
rect 85 15 100 585
rect 50 0 100 15
rect 150 585 200 600
rect 150 15 165 585
rect 185 15 200 585
rect 150 0 200 15
rect 250 585 300 600
rect 350 585 400 600
rect 250 15 265 585
rect 285 15 300 585
rect 350 15 365 585
rect 385 15 400 585
rect 250 0 300 15
rect 350 0 400 15
rect 450 585 500 600
rect 450 15 465 585
rect 485 15 500 585
rect 450 0 500 15
rect 550 585 600 600
rect 550 15 565 585
rect 585 15 600 585
rect 550 0 600 15
rect 650 585 700 600
rect 650 15 665 585
rect 685 15 700 585
rect 650 0 700 15
<< pdiff >>
rect -50 2585 0 2600
rect -50 2015 -35 2585
rect -15 2015 0 2585
rect -50 2000 0 2015
rect 50 2585 100 2600
rect 50 2015 65 2585
rect 85 2015 100 2585
rect 50 2000 100 2015
rect 150 2585 200 2600
rect 150 2015 165 2585
rect 185 2015 200 2585
rect 150 2000 200 2015
rect 250 2585 300 2600
rect 350 2585 400 2600
rect 250 2015 265 2585
rect 285 2015 300 2585
rect 350 2015 365 2585
rect 385 2015 400 2585
rect 250 2000 300 2015
rect 350 2000 400 2015
rect 450 2585 500 2600
rect 450 2015 465 2585
rect 485 2015 500 2585
rect 450 2000 500 2015
rect 550 2585 600 2600
rect 550 2015 565 2585
rect 585 2015 600 2585
rect 550 2000 600 2015
rect 650 2585 700 2600
rect 650 2015 665 2585
rect 685 2015 700 2585
rect 650 2000 700 2015
rect -50 1585 0 1600
rect -50 1015 -35 1585
rect -15 1015 0 1585
rect -50 1000 0 1015
rect 50 1585 100 1600
rect 50 1015 65 1585
rect 85 1015 100 1585
rect 50 1000 100 1015
rect 150 1585 200 1600
rect 150 1015 165 1585
rect 185 1015 200 1585
rect 150 1000 200 1015
rect 250 1585 300 1600
rect 350 1585 400 1600
rect 250 1015 265 1585
rect 285 1015 300 1585
rect 350 1015 365 1585
rect 385 1015 400 1585
rect 250 1000 300 1015
rect 350 1000 400 1015
rect 450 1585 500 1600
rect 450 1015 465 1585
rect 485 1015 500 1585
rect 450 1000 500 1015
rect 550 1585 600 1600
rect 550 1015 565 1585
rect 585 1015 600 1585
rect 550 1000 600 1015
rect 650 1585 700 1600
rect 650 1015 665 1585
rect 685 1015 700 1585
rect 650 1000 700 1015
<< ndiffc >>
rect -35 15 -15 585
rect 65 15 85 585
rect 165 15 185 585
rect 265 15 285 585
rect 365 15 385 585
rect 465 15 485 585
rect 565 15 585 585
rect 665 15 685 585
<< pdiffc >>
rect -35 2015 -15 2585
rect 65 2015 85 2585
rect 165 2015 185 2585
rect 265 2015 285 2585
rect 365 2015 385 2585
rect 465 2015 485 2585
rect 565 2015 585 2585
rect 665 2015 685 2585
rect -35 1015 -15 1585
rect 65 1015 85 1585
rect 165 1015 185 1585
rect 265 1015 285 1585
rect 365 1015 385 1585
rect 465 1015 485 1585
rect 565 1015 585 1585
rect 665 1015 685 1585
<< psubdiff >>
rect 300 585 350 600
rect 300 15 315 585
rect 335 15 350 585
rect 300 0 350 15
<< nsubdiff >>
rect 300 2585 350 2600
rect 300 2015 315 2585
rect 335 2015 350 2585
rect 300 2000 350 2015
rect 300 1585 350 1600
rect 300 1015 315 1585
rect 335 1015 350 1585
rect 300 1000 350 1015
<< psubdiffcont >>
rect 315 15 335 585
<< nsubdiffcont >>
rect 315 2015 335 2585
rect 315 1015 335 1585
<< poly >>
rect 0 2600 50 2620
rect 100 2600 150 2620
rect 200 2600 250 2620
rect 400 2600 450 2620
rect 500 2600 550 2620
rect 600 2600 650 2620
rect 0 1985 50 2000
rect 100 1985 150 2000
rect 200 1985 250 2000
rect 400 1985 450 2000
rect 500 1985 550 2000
rect 600 1985 650 2000
rect 0 1600 50 1620
rect 100 1600 150 1620
rect 200 1600 250 1620
rect 400 1600 450 1620
rect 500 1600 550 1620
rect 600 1600 650 1620
rect 0 985 50 1000
rect 100 985 150 1000
rect 200 985 250 1000
rect 400 985 450 1000
rect 500 985 550 1000
rect 600 985 650 1000
rect 0 600 50 620
rect 100 600 150 615
rect 200 600 250 615
rect 400 600 450 615
rect 500 600 550 615
rect 600 600 650 620
rect 0 -65 50 0
rect 100 -25 150 0
rect 200 -15 250 0
rect 400 -15 450 0
rect 100 -45 115 -25
rect 135 -45 150 -25
rect 100 -60 150 -45
rect 500 -25 550 0
rect 500 -45 515 -25
rect 535 -45 550 -25
rect 500 -60 550 -45
rect 0 -85 15 -65
rect 35 -85 50 -65
rect 0 -100 50 -85
rect 600 -65 650 0
rect 600 -85 615 -65
rect 635 -85 650 -65
rect 600 -100 650 -85
<< polycont >>
rect 115 -45 135 -25
rect 515 -45 535 -25
rect 15 -85 35 -65
rect 615 -85 635 -65
<< locali >>
rect -50 2585 -5 2595
rect -50 2015 -35 2585
rect -15 2015 -5 2585
rect -50 2005 -5 2015
rect 55 2585 95 2595
rect 55 2015 65 2585
rect 85 2015 95 2585
rect 55 2005 95 2015
rect 155 2585 195 2595
rect 155 2015 165 2585
rect 185 2015 195 2585
rect 155 2005 195 2015
rect 255 2585 395 2595
rect 255 2015 265 2585
rect 285 2015 315 2585
rect 335 2015 365 2585
rect 385 2015 395 2585
rect 255 2005 395 2015
rect 455 2585 495 2595
rect 455 2015 465 2585
rect 485 2015 495 2585
rect 455 2005 495 2015
rect 555 2585 595 2595
rect 555 2015 565 2585
rect 585 2015 595 2585
rect 555 2005 595 2015
rect 655 2585 700 2595
rect 655 2015 665 2585
rect 685 2015 700 2585
rect 655 2005 700 2015
rect -50 1585 -5 1595
rect -50 1015 -35 1585
rect -15 1015 -5 1585
rect -50 1005 -5 1015
rect 55 1585 95 1595
rect 55 1015 65 1585
rect 85 1015 95 1585
rect 55 1005 95 1015
rect 155 1585 195 1595
rect 155 1015 165 1585
rect 185 1015 195 1585
rect 155 1005 195 1015
rect 255 1585 395 1595
rect 255 1015 265 1585
rect 285 1015 315 1585
rect 335 1015 365 1585
rect 385 1015 395 1585
rect 255 1005 395 1015
rect 455 1585 495 1595
rect 455 1015 465 1585
rect 485 1015 495 1585
rect 455 1005 495 1015
rect 555 1585 595 1595
rect 555 1015 565 1585
rect 585 1015 595 1585
rect 555 1005 595 1015
rect 655 1585 700 1595
rect 655 1015 665 1585
rect 685 1015 700 1585
rect 655 1005 700 1015
rect -50 585 -5 595
rect -50 15 -35 585
rect -15 15 -5 585
rect -50 5 -5 15
rect 55 585 95 595
rect 55 15 65 585
rect 85 15 95 585
rect 55 5 95 15
rect 155 585 195 595
rect 155 15 165 585
rect 185 15 195 585
rect 155 5 195 15
rect 255 585 395 595
rect 255 15 265 585
rect 285 15 315 585
rect 335 15 365 585
rect 385 15 395 585
rect 255 5 395 15
rect 455 585 495 595
rect 455 15 465 585
rect 485 15 495 585
rect 455 5 495 15
rect 555 585 595 595
rect 555 15 565 585
rect 585 15 595 585
rect 555 5 595 15
rect 655 585 700 595
rect 655 15 665 585
rect 685 15 700 585
rect 655 5 700 15
rect 105 -25 545 -15
rect 105 -45 115 -25
rect 135 -45 515 -25
rect 535 -45 545 -25
rect 105 -55 545 -45
rect 5 -65 45 -55
rect 5 -85 15 -65
rect 35 -75 45 -65
rect 605 -65 645 -55
rect 605 -75 615 -65
rect 35 -85 615 -75
rect 635 -85 645 -65
rect 5 -95 645 -85
<< viali >>
rect 265 2015 285 2585
rect 315 2015 335 2585
rect 365 2015 385 2585
rect 265 1015 285 1585
rect 315 1015 335 1585
rect 365 1015 385 1585
rect 265 15 285 585
rect 315 15 335 585
rect 365 15 385 585
<< metal1 >>
rect -50 2585 700 2600
rect -50 2015 265 2585
rect 285 2015 315 2585
rect 335 2015 365 2585
rect 385 2015 700 2585
rect -50 2000 700 2015
rect -50 1585 700 1600
rect -50 1015 265 1585
rect 285 1015 315 1585
rect 335 1015 365 1585
rect 385 1015 700 1585
rect -50 1000 700 1015
rect -50 585 700 600
rect -50 15 265 585
rect 285 15 315 585
rect 335 15 365 585
rect 385 15 700 585
rect -50 0 700 15
<< end >>
