* SPICE3 file created from inverter.ext - technology: sky130A


* Top level circuit inverter

X0 gnd d ~d gnd sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X1 vdd d ~d vdd sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
.end

